// Generator : SpinalHDL v1.4.3    git head : adf552d8f500e7419fff395b7049228e4bc5de26
// Component : TopLevel
// Git hash  : 772db2e021a60a74f3e57a7af123ee75a269deec


`define UartParityType_defaultEncoding_type [1:0]
`define UartParityType_defaultEncoding_NONE 2'b00
`define UartParityType_defaultEncoding_EVEN 2'b01
`define UartParityType_defaultEncoding_ODD 2'b10

`define UartStopType_defaultEncoding_type [0:0]
`define UartStopType_defaultEncoding_ONE 1'b0
`define UartStopType_defaultEncoding_TWO 1'b1

`define UartCtrlTxState_defaultEncoding_type [2:0]
`define UartCtrlTxState_defaultEncoding_IDLE 3'b000
`define UartCtrlTxState_defaultEncoding_START 3'b001
`define UartCtrlTxState_defaultEncoding_DATA 3'b010
`define UartCtrlTxState_defaultEncoding_PARITY 3'b011
`define UartCtrlTxState_defaultEncoding_STOP 3'b100

`define UartCtrlRxState_defaultEncoding_type [2:0]
`define UartCtrlRxState_defaultEncoding_IDLE 3'b000
`define UartCtrlRxState_defaultEncoding_START 3'b001
`define UartCtrlRxState_defaultEncoding_DATA 3'b010
`define UartCtrlRxState_defaultEncoding_PARITY 3'b011
`define UartCtrlRxState_defaultEncoding_STOP 3'b100

`define machine_enumDefinition_defaultEncoding_type [3:0]
`define machine_enumDefinition_defaultEncoding_machine_BOOT 4'b0000
`define machine_enumDefinition_defaultEncoding_machine_idle 4'b0001
`define machine_enumDefinition_defaultEncoding_machine_k6 4'b0010
`define machine_enumDefinition_defaultEncoding_machine_k5 4'b0011
`define machine_enumDefinition_defaultEncoding_machine_k4 4'b0100
`define machine_enumDefinition_defaultEncoding_machine_k3 4'b0101
`define machine_enumDefinition_defaultEncoding_machine_k2 4'b0110
`define machine_enumDefinition_defaultEncoding_machine_k1 4'b0111
`define machine_enumDefinition_defaultEncoding_machine_reserved 4'b1000
`define machine_enumDefinition_defaultEncoding_machine_special 4'b1001


module TopLevel (
  input               KEY_Fn,
  input               CLK_50,
  input      [20:0]   COL,
  output     [5:0]    LED_A,
  output     [5:0]    ROW,
  output     [34:0]   LED_K,
  output              TXD,
  output              LED_R6,
   inout              PS2_CLK,
   inout              PS2_DAT,
  output              flash_dclk,
  output              flash_sce,
  output              flash_sdo,
  input               flash_data0
);
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire       [2:0]    _zz_8;
  wire       `UartStopType_defaultEncoding_type _zz_9;
  wire       `UartParityType_defaultEncoding_type _zz_10;
  wire       [19:0]   _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire                _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire                _zz_152;
  wire                _zz_153;
  wire                _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire                _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire                _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire                _zz_170;
  wire                _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire                _zz_174;
  wire                _zz_175;
  wire                _zz_176;
  wire                _zz_177;
  wire                _zz_178;
  wire                _zz_179;
  wire                _zz_180;
  wire                _zz_181;
  wire                _zz_182;
  wire                _zz_183;
  wire                _zz_184;
  wire                _zz_185;
  wire                _zz_186;
  wire                _zz_187;
  wire                _zz_188;
  wire                _zz_189;
  wire                _zz_190;
  wire                _zz_191;
  wire                _zz_192;
  wire                _zz_193;
  wire                _zz_194;
  wire                _zz_195;
  wire                _zz_196;
  wire                _zz_197;
  wire                _zz_198;
  wire                _zz_199;
  wire                _zz_200;
  wire                _zz_201;
  wire                _zz_202;
  wire                _zz_203;
  wire                _zz_204;
  wire                _zz_205;
  wire                _zz_206;
  wire                pll100_c0;
  wire                pll100_locked;
  wire                rstCtrl_io_globalReset;
  wire                bufferCC_3_io_dataOut;
  wire                core_uart_txd;
  wire       [5:0]    core_io_row;
  wire       [34:0]   core_io_col;
  wire                core_flash_dclk;
  wire                core_flash_sce;
  wire                core_flash_sdo;
  wire       [5:0]    clk50Area_keyMatrix_ROW;
  wire                clk50Area_keyMatrix_scanIdx_valid;
  wire       [7:0]    clk50Area_keyMatrix_scanIdx_payload;
  wire                clk50Area_keyMatrix_keyStatus_0_valid;
  wire                clk50Area_keyMatrix_keyStatus_0_payload;
  wire                clk50Area_keyMatrix_keyStatus_1_valid;
  wire                clk50Area_keyMatrix_keyStatus_1_payload;
  wire                clk50Area_keyMatrix_keyStatus_2_valid;
  wire                clk50Area_keyMatrix_keyStatus_2_payload;
  wire                clk50Area_keyMatrix_keyStatus_3_valid;
  wire                clk50Area_keyMatrix_keyStatus_3_payload;
  wire                clk50Area_keyMatrix_keyStatus_4_valid;
  wire                clk50Area_keyMatrix_keyStatus_4_payload;
  wire                clk50Area_keyMatrix_keyStatus_5_valid;
  wire                clk50Area_keyMatrix_keyStatus_5_payload;
  wire                clk50Area_keyMatrix_keyStatus_6_valid;
  wire                clk50Area_keyMatrix_keyStatus_6_payload;
  wire                clk50Area_keyMatrix_keyStatus_7_valid;
  wire                clk50Area_keyMatrix_keyStatus_7_payload;
  wire                clk50Area_keyMatrix_keyStatus_8_valid;
  wire                clk50Area_keyMatrix_keyStatus_8_payload;
  wire                clk50Area_keyMatrix_keyStatus_9_valid;
  wire                clk50Area_keyMatrix_keyStatus_9_payload;
  wire                clk50Area_keyMatrix_keyStatus_10_valid;
  wire                clk50Area_keyMatrix_keyStatus_10_payload;
  wire                clk50Area_keyMatrix_keyStatus_11_valid;
  wire                clk50Area_keyMatrix_keyStatus_11_payload;
  wire                clk50Area_keyMatrix_keyStatus_12_valid;
  wire                clk50Area_keyMatrix_keyStatus_12_payload;
  wire                clk50Area_keyMatrix_keyStatus_13_valid;
  wire                clk50Area_keyMatrix_keyStatus_13_payload;
  wire                clk50Area_keyMatrix_keyStatus_14_valid;
  wire                clk50Area_keyMatrix_keyStatus_14_payload;
  wire                clk50Area_keyMatrix_keyStatus_15_valid;
  wire                clk50Area_keyMatrix_keyStatus_15_payload;
  wire                clk50Area_keyMatrix_keyStatus_16_valid;
  wire                clk50Area_keyMatrix_keyStatus_16_payload;
  wire                clk50Area_keyMatrix_keyStatus_17_valid;
  wire                clk50Area_keyMatrix_keyStatus_17_payload;
  wire                clk50Area_keyMatrix_keyStatus_18_valid;
  wire                clk50Area_keyMatrix_keyStatus_18_payload;
  wire                clk50Area_keyMatrix_keyStatus_19_valid;
  wire                clk50Area_keyMatrix_keyStatus_19_payload;
  wire                clk50Area_keyMatrix_keyStatus_20_valid;
  wire                clk50Area_keyMatrix_keyStatus_20_payload;
  wire                clk50Area_keyMatrix_keyStatus_21_valid;
  wire                clk50Area_keyMatrix_keyStatus_21_payload;
  wire                clk50Area_keyMatrix_keyStatus_22_valid;
  wire                clk50Area_keyMatrix_keyStatus_22_payload;
  wire                clk50Area_keyMatrix_keyStatus_23_valid;
  wire                clk50Area_keyMatrix_keyStatus_23_payload;
  wire                clk50Area_keyMatrix_keyStatus_24_valid;
  wire                clk50Area_keyMatrix_keyStatus_24_payload;
  wire                clk50Area_keyMatrix_keyStatus_25_valid;
  wire                clk50Area_keyMatrix_keyStatus_25_payload;
  wire                clk50Area_keyMatrix_keyStatus_26_valid;
  wire                clk50Area_keyMatrix_keyStatus_26_payload;
  wire                clk50Area_keyMatrix_keyStatus_27_valid;
  wire                clk50Area_keyMatrix_keyStatus_27_payload;
  wire                clk50Area_keyMatrix_keyStatus_28_valid;
  wire                clk50Area_keyMatrix_keyStatus_28_payload;
  wire                clk50Area_keyMatrix_keyStatus_29_valid;
  wire                clk50Area_keyMatrix_keyStatus_29_payload;
  wire                clk50Area_keyMatrix_keyStatus_30_valid;
  wire                clk50Area_keyMatrix_keyStatus_30_payload;
  wire                clk50Area_keyMatrix_keyStatus_31_valid;
  wire                clk50Area_keyMatrix_keyStatus_31_payload;
  wire                clk50Area_keyMatrix_keyStatus_32_valid;
  wire                clk50Area_keyMatrix_keyStatus_32_payload;
  wire                clk50Area_keyMatrix_keyStatus_33_valid;
  wire                clk50Area_keyMatrix_keyStatus_33_payload;
  wire                clk50Area_keyMatrix_keyStatus_34_valid;
  wire                clk50Area_keyMatrix_keyStatus_34_payload;
  wire                clk50Area_keyMatrix_keyStatus_35_valid;
  wire                clk50Area_keyMatrix_keyStatus_35_payload;
  wire                clk50Area_keyMatrix_keyStatus_36_valid;
  wire                clk50Area_keyMatrix_keyStatus_36_payload;
  wire                clk50Area_keyMatrix_keyStatus_37_valid;
  wire                clk50Area_keyMatrix_keyStatus_37_payload;
  wire                clk50Area_keyMatrix_keyStatus_38_valid;
  wire                clk50Area_keyMatrix_keyStatus_38_payload;
  wire                clk50Area_keyMatrix_keyStatus_39_valid;
  wire                clk50Area_keyMatrix_keyStatus_39_payload;
  wire                clk50Area_keyMatrix_keyStatus_40_valid;
  wire                clk50Area_keyMatrix_keyStatus_40_payload;
  wire                clk50Area_keyMatrix_keyStatus_41_valid;
  wire                clk50Area_keyMatrix_keyStatus_41_payload;
  wire                clk50Area_keyMatrix_keyStatus_42_valid;
  wire                clk50Area_keyMatrix_keyStatus_42_payload;
  wire                clk50Area_keyMatrix_keyStatus_43_valid;
  wire                clk50Area_keyMatrix_keyStatus_43_payload;
  wire                clk50Area_keyMatrix_keyStatus_44_valid;
  wire                clk50Area_keyMatrix_keyStatus_44_payload;
  wire                clk50Area_keyMatrix_keyStatus_45_valid;
  wire                clk50Area_keyMatrix_keyStatus_45_payload;
  wire                clk50Area_keyMatrix_keyStatus_46_valid;
  wire                clk50Area_keyMatrix_keyStatus_46_payload;
  wire                clk50Area_keyMatrix_keyStatus_47_valid;
  wire                clk50Area_keyMatrix_keyStatus_47_payload;
  wire                clk50Area_keyMatrix_keyStatus_48_valid;
  wire                clk50Area_keyMatrix_keyStatus_48_payload;
  wire                clk50Area_keyMatrix_keyStatus_49_valid;
  wire                clk50Area_keyMatrix_keyStatus_49_payload;
  wire                clk50Area_keyMatrix_keyStatus_50_valid;
  wire                clk50Area_keyMatrix_keyStatus_50_payload;
  wire                clk50Area_keyMatrix_keyStatus_51_valid;
  wire                clk50Area_keyMatrix_keyStatus_51_payload;
  wire                clk50Area_keyMatrix_keyStatus_52_valid;
  wire                clk50Area_keyMatrix_keyStatus_52_payload;
  wire                clk50Area_keyMatrix_keyStatus_53_valid;
  wire                clk50Area_keyMatrix_keyStatus_53_payload;
  wire                clk50Area_keyMatrix_keyStatus_54_valid;
  wire                clk50Area_keyMatrix_keyStatus_54_payload;
  wire                clk50Area_keyMatrix_keyStatus_55_valid;
  wire                clk50Area_keyMatrix_keyStatus_55_payload;
  wire                clk50Area_keyMatrix_keyStatus_56_valid;
  wire                clk50Area_keyMatrix_keyStatus_56_payload;
  wire                clk50Area_keyMatrix_keyStatus_57_valid;
  wire                clk50Area_keyMatrix_keyStatus_57_payload;
  wire                clk50Area_keyMatrix_keyStatus_58_valid;
  wire                clk50Area_keyMatrix_keyStatus_58_payload;
  wire                clk50Area_keyMatrix_keyStatus_59_valid;
  wire                clk50Area_keyMatrix_keyStatus_59_payload;
  wire                clk50Area_keyMatrix_keyStatus_60_valid;
  wire                clk50Area_keyMatrix_keyStatus_60_payload;
  wire                clk50Area_keyMatrix_keyStatus_61_valid;
  wire                clk50Area_keyMatrix_keyStatus_61_payload;
  wire                clk50Area_keyMatrix_keyStatus_62_valid;
  wire                clk50Area_keyMatrix_keyStatus_62_payload;
  wire                clk50Area_keyMatrix_keyStatus_63_valid;
  wire                clk50Area_keyMatrix_keyStatus_63_payload;
  wire                clk50Area_keyMatrix_keyStatus_64_valid;
  wire                clk50Area_keyMatrix_keyStatus_64_payload;
  wire                clk50Area_keyMatrix_keyStatus_65_valid;
  wire                clk50Area_keyMatrix_keyStatus_65_payload;
  wire                clk50Area_keyMatrix_keyStatus_66_valid;
  wire                clk50Area_keyMatrix_keyStatus_66_payload;
  wire                clk50Area_keyMatrix_keyStatus_67_valid;
  wire                clk50Area_keyMatrix_keyStatus_67_payload;
  wire                clk50Area_keyMatrix_keyStatus_68_valid;
  wire                clk50Area_keyMatrix_keyStatus_68_payload;
  wire                clk50Area_keyMatrix_keyStatus_69_valid;
  wire                clk50Area_keyMatrix_keyStatus_69_payload;
  wire                clk50Area_keyMatrix_keyStatus_70_valid;
  wire                clk50Area_keyMatrix_keyStatus_70_payload;
  wire                clk50Area_keyMatrix_keyStatus_71_valid;
  wire                clk50Area_keyMatrix_keyStatus_71_payload;
  wire                clk50Area_keyMatrix_keyStatus_72_valid;
  wire                clk50Area_keyMatrix_keyStatus_72_payload;
  wire                clk50Area_keyMatrix_keyStatus_73_valid;
  wire                clk50Area_keyMatrix_keyStatus_73_payload;
  wire                clk50Area_keyMatrix_keyStatus_74_valid;
  wire                clk50Area_keyMatrix_keyStatus_74_payload;
  wire                clk50Area_keyMatrix_keyStatus_75_valid;
  wire                clk50Area_keyMatrix_keyStatus_75_payload;
  wire                clk50Area_keyMatrix_keyStatus_76_valid;
  wire                clk50Area_keyMatrix_keyStatus_76_payload;
  wire                clk50Area_keyMatrix_keyStatus_77_valid;
  wire                clk50Area_keyMatrix_keyStatus_77_payload;
  wire                clk50Area_keyMatrix_keyStatus_78_valid;
  wire                clk50Area_keyMatrix_keyStatus_78_payload;
  wire                clk50Area_keyMatrix_keyStatus_79_valid;
  wire                clk50Area_keyMatrix_keyStatus_79_payload;
  wire                clk50Area_keyMatrix_keyStatus_80_valid;
  wire                clk50Area_keyMatrix_keyStatus_80_payload;
  wire                clk50Area_keyMatrix_keyStatus_81_valid;
  wire                clk50Area_keyMatrix_keyStatus_81_payload;
  wire                clk50Area_keyMatrix_keyStatus_82_valid;
  wire                clk50Area_keyMatrix_keyStatus_82_payload;
  wire                clk50Area_keyMatrix_keyStatus_83_valid;
  wire                clk50Area_keyMatrix_keyStatus_83_payload;
  wire                clk50Area_keyMatrix_keyStatus_84_valid;
  wire                clk50Area_keyMatrix_keyStatus_84_payload;
  wire                clk50Area_keyMatrix_keyStatus_85_valid;
  wire                clk50Area_keyMatrix_keyStatus_85_payload;
  wire                clk50Area_keyMatrix_keyStatus_86_valid;
  wire                clk50Area_keyMatrix_keyStatus_86_payload;
  wire                clk50Area_keyMatrix_keyStatus_87_valid;
  wire                clk50Area_keyMatrix_keyStatus_87_payload;
  wire                clk50Area_keyMatrix_keyStatus_88_valid;
  wire                clk50Area_keyMatrix_keyStatus_88_payload;
  wire                clk50Area_keyMatrix_keyStatus_89_valid;
  wire                clk50Area_keyMatrix_keyStatus_89_payload;
  wire                clk50Area_keyMatrix_keyStatus_90_valid;
  wire                clk50Area_keyMatrix_keyStatus_90_payload;
  wire                clk50Area_keyMatrix_keyStatus_91_valid;
  wire                clk50Area_keyMatrix_keyStatus_91_payload;
  wire                clk50Area_keyMatrix_keyStatus_92_valid;
  wire                clk50Area_keyMatrix_keyStatus_92_payload;
  wire                clk50Area_keyMatrix_keyStatus_93_valid;
  wire                clk50Area_keyMatrix_keyStatus_93_payload;
  wire                clk50Area_keyMatrix_keyStatus_94_valid;
  wire                clk50Area_keyMatrix_keyStatus_94_payload;
  wire                clk50Area_keyMatrix_keyStatus_95_valid;
  wire                clk50Area_keyMatrix_keyStatus_95_payload;
  wire                clk50Area_keyMatrix_keyStatus_96_valid;
  wire                clk50Area_keyMatrix_keyStatus_96_payload;
  wire                clk50Area_keyMatrix_keyStatus_97_valid;
  wire                clk50Area_keyMatrix_keyStatus_97_payload;
  wire                clk50Area_keyMatrix_keyStatus_98_valid;
  wire                clk50Area_keyMatrix_keyStatus_98_payload;
  wire                clk50Area_keyMatrix_keyStatus_99_valid;
  wire                clk50Area_keyMatrix_keyStatus_99_payload;
  wire                clk50Area_keyMatrix_keyStatus_100_valid;
  wire                clk50Area_keyMatrix_keyStatus_100_payload;
  wire                clk50Area_keyMatrix_keyStatus_101_valid;
  wire                clk50Area_keyMatrix_keyStatus_101_payload;
  wire                clk50Area_keyMatrix_keyStatus_102_valid;
  wire                clk50Area_keyMatrix_keyStatus_102_payload;
  wire                uartCtrl_2_io_write_ready;
  wire                uartCtrl_2_io_read_valid;
  wire       [7:0]    uartCtrl_2_io_read_payload;
  wire                uartCtrl_2_io_uart_txd;
  wire                uartCtrl_2_io_readError;
  wire                uartCtrl_2_io_readBreak;
  wire                clk50Area_hid_TXD;
  reg                 _zz_1;
  wire                _zz_2;
  reg        [7:0]    clk50Area_keyMatrix_scanIdx_payload_regNextWhen;
  reg                 _zz_3;

  pll pll100 (
    .inclk0    (CLK_50         ), //i
    .c0        (pll100_c0      ), //o
    .locked    (pll100_locked  )  //o
  );
  ResetController rstCtrl (
    .io_clock            (CLK_50                  ), //i
    .io_externalReset    (_zz_4                   ), //i
    .io_globalReset      (rstCtrl_io_globalReset  )  //o
  );
  BufferCC_2 bufferCC_3 (
    .io_dataIn     (_zz_5                  ), //i
    .io_dataOut    (bufferCC_3_io_dataOut  ), //o
    .CLK_50        (CLK_50                 ), //i
    ._zz_1         (_zz_2                  )  //i
  );
  kbd104 core (
    .clk_clk          (pll100_c0               ), //i
    .reset_reset_n    (_zz_6                   ), //i
    .uart_txd         (core_uart_txd           ), //o
    .uart_rxd         (uartCtrl_2_io_uart_txd  ), //i
    .io_row           (core_io_row[5:0]        ), //o
    .io_col           (core_io_col[34:0]       ), //o
    .flash_dclk       (core_flash_dclk         ), //o
    .flash_sce        (core_flash_sce          ), //o
    .flash_sdo        (core_flash_sdo          ), //o
    .flash_data0      (flash_data0             )  //i
  );
  KeyMatrix clk50Area_keyMatrix (
    .enabled                  (_zz_7                                      ), //i
    .COL                      (COL[20:0]                                  ), //i
    .ROW                      (clk50Area_keyMatrix_ROW[5:0]               ), //o
    .scanIdx_valid            (clk50Area_keyMatrix_scanIdx_valid          ), //o
    .scanIdx_payload          (clk50Area_keyMatrix_scanIdx_payload[7:0]   ), //o
    .keyStatus_0_valid        (clk50Area_keyMatrix_keyStatus_0_valid      ), //o
    .keyStatus_0_payload      (clk50Area_keyMatrix_keyStatus_0_payload    ), //o
    .keyStatus_1_valid        (clk50Area_keyMatrix_keyStatus_1_valid      ), //o
    .keyStatus_1_payload      (clk50Area_keyMatrix_keyStatus_1_payload    ), //o
    .keyStatus_2_valid        (clk50Area_keyMatrix_keyStatus_2_valid      ), //o
    .keyStatus_2_payload      (clk50Area_keyMatrix_keyStatus_2_payload    ), //o
    .keyStatus_3_valid        (clk50Area_keyMatrix_keyStatus_3_valid      ), //o
    .keyStatus_3_payload      (clk50Area_keyMatrix_keyStatus_3_payload    ), //o
    .keyStatus_4_valid        (clk50Area_keyMatrix_keyStatus_4_valid      ), //o
    .keyStatus_4_payload      (clk50Area_keyMatrix_keyStatus_4_payload    ), //o
    .keyStatus_5_valid        (clk50Area_keyMatrix_keyStatus_5_valid      ), //o
    .keyStatus_5_payload      (clk50Area_keyMatrix_keyStatus_5_payload    ), //o
    .keyStatus_6_valid        (clk50Area_keyMatrix_keyStatus_6_valid      ), //o
    .keyStatus_6_payload      (clk50Area_keyMatrix_keyStatus_6_payload    ), //o
    .keyStatus_7_valid        (clk50Area_keyMatrix_keyStatus_7_valid      ), //o
    .keyStatus_7_payload      (clk50Area_keyMatrix_keyStatus_7_payload    ), //o
    .keyStatus_8_valid        (clk50Area_keyMatrix_keyStatus_8_valid      ), //o
    .keyStatus_8_payload      (clk50Area_keyMatrix_keyStatus_8_payload    ), //o
    .keyStatus_9_valid        (clk50Area_keyMatrix_keyStatus_9_valid      ), //o
    .keyStatus_9_payload      (clk50Area_keyMatrix_keyStatus_9_payload    ), //o
    .keyStatus_10_valid       (clk50Area_keyMatrix_keyStatus_10_valid     ), //o
    .keyStatus_10_payload     (clk50Area_keyMatrix_keyStatus_10_payload   ), //o
    .keyStatus_11_valid       (clk50Area_keyMatrix_keyStatus_11_valid     ), //o
    .keyStatus_11_payload     (clk50Area_keyMatrix_keyStatus_11_payload   ), //o
    .keyStatus_12_valid       (clk50Area_keyMatrix_keyStatus_12_valid     ), //o
    .keyStatus_12_payload     (clk50Area_keyMatrix_keyStatus_12_payload   ), //o
    .keyStatus_13_valid       (clk50Area_keyMatrix_keyStatus_13_valid     ), //o
    .keyStatus_13_payload     (clk50Area_keyMatrix_keyStatus_13_payload   ), //o
    .keyStatus_14_valid       (clk50Area_keyMatrix_keyStatus_14_valid     ), //o
    .keyStatus_14_payload     (clk50Area_keyMatrix_keyStatus_14_payload   ), //o
    .keyStatus_15_valid       (clk50Area_keyMatrix_keyStatus_15_valid     ), //o
    .keyStatus_15_payload     (clk50Area_keyMatrix_keyStatus_15_payload   ), //o
    .keyStatus_16_valid       (clk50Area_keyMatrix_keyStatus_16_valid     ), //o
    .keyStatus_16_payload     (clk50Area_keyMatrix_keyStatus_16_payload   ), //o
    .keyStatus_17_valid       (clk50Area_keyMatrix_keyStatus_17_valid     ), //o
    .keyStatus_17_payload     (clk50Area_keyMatrix_keyStatus_17_payload   ), //o
    .keyStatus_18_valid       (clk50Area_keyMatrix_keyStatus_18_valid     ), //o
    .keyStatus_18_payload     (clk50Area_keyMatrix_keyStatus_18_payload   ), //o
    .keyStatus_19_valid       (clk50Area_keyMatrix_keyStatus_19_valid     ), //o
    .keyStatus_19_payload     (clk50Area_keyMatrix_keyStatus_19_payload   ), //o
    .keyStatus_20_valid       (clk50Area_keyMatrix_keyStatus_20_valid     ), //o
    .keyStatus_20_payload     (clk50Area_keyMatrix_keyStatus_20_payload   ), //o
    .keyStatus_21_valid       (clk50Area_keyMatrix_keyStatus_21_valid     ), //o
    .keyStatus_21_payload     (clk50Area_keyMatrix_keyStatus_21_payload   ), //o
    .keyStatus_22_valid       (clk50Area_keyMatrix_keyStatus_22_valid     ), //o
    .keyStatus_22_payload     (clk50Area_keyMatrix_keyStatus_22_payload   ), //o
    .keyStatus_23_valid       (clk50Area_keyMatrix_keyStatus_23_valid     ), //o
    .keyStatus_23_payload     (clk50Area_keyMatrix_keyStatus_23_payload   ), //o
    .keyStatus_24_valid       (clk50Area_keyMatrix_keyStatus_24_valid     ), //o
    .keyStatus_24_payload     (clk50Area_keyMatrix_keyStatus_24_payload   ), //o
    .keyStatus_25_valid       (clk50Area_keyMatrix_keyStatus_25_valid     ), //o
    .keyStatus_25_payload     (clk50Area_keyMatrix_keyStatus_25_payload   ), //o
    .keyStatus_26_valid       (clk50Area_keyMatrix_keyStatus_26_valid     ), //o
    .keyStatus_26_payload     (clk50Area_keyMatrix_keyStatus_26_payload   ), //o
    .keyStatus_27_valid       (clk50Area_keyMatrix_keyStatus_27_valid     ), //o
    .keyStatus_27_payload     (clk50Area_keyMatrix_keyStatus_27_payload   ), //o
    .keyStatus_28_valid       (clk50Area_keyMatrix_keyStatus_28_valid     ), //o
    .keyStatus_28_payload     (clk50Area_keyMatrix_keyStatus_28_payload   ), //o
    .keyStatus_29_valid       (clk50Area_keyMatrix_keyStatus_29_valid     ), //o
    .keyStatus_29_payload     (clk50Area_keyMatrix_keyStatus_29_payload   ), //o
    .keyStatus_30_valid       (clk50Area_keyMatrix_keyStatus_30_valid     ), //o
    .keyStatus_30_payload     (clk50Area_keyMatrix_keyStatus_30_payload   ), //o
    .keyStatus_31_valid       (clk50Area_keyMatrix_keyStatus_31_valid     ), //o
    .keyStatus_31_payload     (clk50Area_keyMatrix_keyStatus_31_payload   ), //o
    .keyStatus_32_valid       (clk50Area_keyMatrix_keyStatus_32_valid     ), //o
    .keyStatus_32_payload     (clk50Area_keyMatrix_keyStatus_32_payload   ), //o
    .keyStatus_33_valid       (clk50Area_keyMatrix_keyStatus_33_valid     ), //o
    .keyStatus_33_payload     (clk50Area_keyMatrix_keyStatus_33_payload   ), //o
    .keyStatus_34_valid       (clk50Area_keyMatrix_keyStatus_34_valid     ), //o
    .keyStatus_34_payload     (clk50Area_keyMatrix_keyStatus_34_payload   ), //o
    .keyStatus_35_valid       (clk50Area_keyMatrix_keyStatus_35_valid     ), //o
    .keyStatus_35_payload     (clk50Area_keyMatrix_keyStatus_35_payload   ), //o
    .keyStatus_36_valid       (clk50Area_keyMatrix_keyStatus_36_valid     ), //o
    .keyStatus_36_payload     (clk50Area_keyMatrix_keyStatus_36_payload   ), //o
    .keyStatus_37_valid       (clk50Area_keyMatrix_keyStatus_37_valid     ), //o
    .keyStatus_37_payload     (clk50Area_keyMatrix_keyStatus_37_payload   ), //o
    .keyStatus_38_valid       (clk50Area_keyMatrix_keyStatus_38_valid     ), //o
    .keyStatus_38_payload     (clk50Area_keyMatrix_keyStatus_38_payload   ), //o
    .keyStatus_39_valid       (clk50Area_keyMatrix_keyStatus_39_valid     ), //o
    .keyStatus_39_payload     (clk50Area_keyMatrix_keyStatus_39_payload   ), //o
    .keyStatus_40_valid       (clk50Area_keyMatrix_keyStatus_40_valid     ), //o
    .keyStatus_40_payload     (clk50Area_keyMatrix_keyStatus_40_payload   ), //o
    .keyStatus_41_valid       (clk50Area_keyMatrix_keyStatus_41_valid     ), //o
    .keyStatus_41_payload     (clk50Area_keyMatrix_keyStatus_41_payload   ), //o
    .keyStatus_42_valid       (clk50Area_keyMatrix_keyStatus_42_valid     ), //o
    .keyStatus_42_payload     (clk50Area_keyMatrix_keyStatus_42_payload   ), //o
    .keyStatus_43_valid       (clk50Area_keyMatrix_keyStatus_43_valid     ), //o
    .keyStatus_43_payload     (clk50Area_keyMatrix_keyStatus_43_payload   ), //o
    .keyStatus_44_valid       (clk50Area_keyMatrix_keyStatus_44_valid     ), //o
    .keyStatus_44_payload     (clk50Area_keyMatrix_keyStatus_44_payload   ), //o
    .keyStatus_45_valid       (clk50Area_keyMatrix_keyStatus_45_valid     ), //o
    .keyStatus_45_payload     (clk50Area_keyMatrix_keyStatus_45_payload   ), //o
    .keyStatus_46_valid       (clk50Area_keyMatrix_keyStatus_46_valid     ), //o
    .keyStatus_46_payload     (clk50Area_keyMatrix_keyStatus_46_payload   ), //o
    .keyStatus_47_valid       (clk50Area_keyMatrix_keyStatus_47_valid     ), //o
    .keyStatus_47_payload     (clk50Area_keyMatrix_keyStatus_47_payload   ), //o
    .keyStatus_48_valid       (clk50Area_keyMatrix_keyStatus_48_valid     ), //o
    .keyStatus_48_payload     (clk50Area_keyMatrix_keyStatus_48_payload   ), //o
    .keyStatus_49_valid       (clk50Area_keyMatrix_keyStatus_49_valid     ), //o
    .keyStatus_49_payload     (clk50Area_keyMatrix_keyStatus_49_payload   ), //o
    .keyStatus_50_valid       (clk50Area_keyMatrix_keyStatus_50_valid     ), //o
    .keyStatus_50_payload     (clk50Area_keyMatrix_keyStatus_50_payload   ), //o
    .keyStatus_51_valid       (clk50Area_keyMatrix_keyStatus_51_valid     ), //o
    .keyStatus_51_payload     (clk50Area_keyMatrix_keyStatus_51_payload   ), //o
    .keyStatus_52_valid       (clk50Area_keyMatrix_keyStatus_52_valid     ), //o
    .keyStatus_52_payload     (clk50Area_keyMatrix_keyStatus_52_payload   ), //o
    .keyStatus_53_valid       (clk50Area_keyMatrix_keyStatus_53_valid     ), //o
    .keyStatus_53_payload     (clk50Area_keyMatrix_keyStatus_53_payload   ), //o
    .keyStatus_54_valid       (clk50Area_keyMatrix_keyStatus_54_valid     ), //o
    .keyStatus_54_payload     (clk50Area_keyMatrix_keyStatus_54_payload   ), //o
    .keyStatus_55_valid       (clk50Area_keyMatrix_keyStatus_55_valid     ), //o
    .keyStatus_55_payload     (clk50Area_keyMatrix_keyStatus_55_payload   ), //o
    .keyStatus_56_valid       (clk50Area_keyMatrix_keyStatus_56_valid     ), //o
    .keyStatus_56_payload     (clk50Area_keyMatrix_keyStatus_56_payload   ), //o
    .keyStatus_57_valid       (clk50Area_keyMatrix_keyStatus_57_valid     ), //o
    .keyStatus_57_payload     (clk50Area_keyMatrix_keyStatus_57_payload   ), //o
    .keyStatus_58_valid       (clk50Area_keyMatrix_keyStatus_58_valid     ), //o
    .keyStatus_58_payload     (clk50Area_keyMatrix_keyStatus_58_payload   ), //o
    .keyStatus_59_valid       (clk50Area_keyMatrix_keyStatus_59_valid     ), //o
    .keyStatus_59_payload     (clk50Area_keyMatrix_keyStatus_59_payload   ), //o
    .keyStatus_60_valid       (clk50Area_keyMatrix_keyStatus_60_valid     ), //o
    .keyStatus_60_payload     (clk50Area_keyMatrix_keyStatus_60_payload   ), //o
    .keyStatus_61_valid       (clk50Area_keyMatrix_keyStatus_61_valid     ), //o
    .keyStatus_61_payload     (clk50Area_keyMatrix_keyStatus_61_payload   ), //o
    .keyStatus_62_valid       (clk50Area_keyMatrix_keyStatus_62_valid     ), //o
    .keyStatus_62_payload     (clk50Area_keyMatrix_keyStatus_62_payload   ), //o
    .keyStatus_63_valid       (clk50Area_keyMatrix_keyStatus_63_valid     ), //o
    .keyStatus_63_payload     (clk50Area_keyMatrix_keyStatus_63_payload   ), //o
    .keyStatus_64_valid       (clk50Area_keyMatrix_keyStatus_64_valid     ), //o
    .keyStatus_64_payload     (clk50Area_keyMatrix_keyStatus_64_payload   ), //o
    .keyStatus_65_valid       (clk50Area_keyMatrix_keyStatus_65_valid     ), //o
    .keyStatus_65_payload     (clk50Area_keyMatrix_keyStatus_65_payload   ), //o
    .keyStatus_66_valid       (clk50Area_keyMatrix_keyStatus_66_valid     ), //o
    .keyStatus_66_payload     (clk50Area_keyMatrix_keyStatus_66_payload   ), //o
    .keyStatus_67_valid       (clk50Area_keyMatrix_keyStatus_67_valid     ), //o
    .keyStatus_67_payload     (clk50Area_keyMatrix_keyStatus_67_payload   ), //o
    .keyStatus_68_valid       (clk50Area_keyMatrix_keyStatus_68_valid     ), //o
    .keyStatus_68_payload     (clk50Area_keyMatrix_keyStatus_68_payload   ), //o
    .keyStatus_69_valid       (clk50Area_keyMatrix_keyStatus_69_valid     ), //o
    .keyStatus_69_payload     (clk50Area_keyMatrix_keyStatus_69_payload   ), //o
    .keyStatus_70_valid       (clk50Area_keyMatrix_keyStatus_70_valid     ), //o
    .keyStatus_70_payload     (clk50Area_keyMatrix_keyStatus_70_payload   ), //o
    .keyStatus_71_valid       (clk50Area_keyMatrix_keyStatus_71_valid     ), //o
    .keyStatus_71_payload     (clk50Area_keyMatrix_keyStatus_71_payload   ), //o
    .keyStatus_72_valid       (clk50Area_keyMatrix_keyStatus_72_valid     ), //o
    .keyStatus_72_payload     (clk50Area_keyMatrix_keyStatus_72_payload   ), //o
    .keyStatus_73_valid       (clk50Area_keyMatrix_keyStatus_73_valid     ), //o
    .keyStatus_73_payload     (clk50Area_keyMatrix_keyStatus_73_payload   ), //o
    .keyStatus_74_valid       (clk50Area_keyMatrix_keyStatus_74_valid     ), //o
    .keyStatus_74_payload     (clk50Area_keyMatrix_keyStatus_74_payload   ), //o
    .keyStatus_75_valid       (clk50Area_keyMatrix_keyStatus_75_valid     ), //o
    .keyStatus_75_payload     (clk50Area_keyMatrix_keyStatus_75_payload   ), //o
    .keyStatus_76_valid       (clk50Area_keyMatrix_keyStatus_76_valid     ), //o
    .keyStatus_76_payload     (clk50Area_keyMatrix_keyStatus_76_payload   ), //o
    .keyStatus_77_valid       (clk50Area_keyMatrix_keyStatus_77_valid     ), //o
    .keyStatus_77_payload     (clk50Area_keyMatrix_keyStatus_77_payload   ), //o
    .keyStatus_78_valid       (clk50Area_keyMatrix_keyStatus_78_valid     ), //o
    .keyStatus_78_payload     (clk50Area_keyMatrix_keyStatus_78_payload   ), //o
    .keyStatus_79_valid       (clk50Area_keyMatrix_keyStatus_79_valid     ), //o
    .keyStatus_79_payload     (clk50Area_keyMatrix_keyStatus_79_payload   ), //o
    .keyStatus_80_valid       (clk50Area_keyMatrix_keyStatus_80_valid     ), //o
    .keyStatus_80_payload     (clk50Area_keyMatrix_keyStatus_80_payload   ), //o
    .keyStatus_81_valid       (clk50Area_keyMatrix_keyStatus_81_valid     ), //o
    .keyStatus_81_payload     (clk50Area_keyMatrix_keyStatus_81_payload   ), //o
    .keyStatus_82_valid       (clk50Area_keyMatrix_keyStatus_82_valid     ), //o
    .keyStatus_82_payload     (clk50Area_keyMatrix_keyStatus_82_payload   ), //o
    .keyStatus_83_valid       (clk50Area_keyMatrix_keyStatus_83_valid     ), //o
    .keyStatus_83_payload     (clk50Area_keyMatrix_keyStatus_83_payload   ), //o
    .keyStatus_84_valid       (clk50Area_keyMatrix_keyStatus_84_valid     ), //o
    .keyStatus_84_payload     (clk50Area_keyMatrix_keyStatus_84_payload   ), //o
    .keyStatus_85_valid       (clk50Area_keyMatrix_keyStatus_85_valid     ), //o
    .keyStatus_85_payload     (clk50Area_keyMatrix_keyStatus_85_payload   ), //o
    .keyStatus_86_valid       (clk50Area_keyMatrix_keyStatus_86_valid     ), //o
    .keyStatus_86_payload     (clk50Area_keyMatrix_keyStatus_86_payload   ), //o
    .keyStatus_87_valid       (clk50Area_keyMatrix_keyStatus_87_valid     ), //o
    .keyStatus_87_payload     (clk50Area_keyMatrix_keyStatus_87_payload   ), //o
    .keyStatus_88_valid       (clk50Area_keyMatrix_keyStatus_88_valid     ), //o
    .keyStatus_88_payload     (clk50Area_keyMatrix_keyStatus_88_payload   ), //o
    .keyStatus_89_valid       (clk50Area_keyMatrix_keyStatus_89_valid     ), //o
    .keyStatus_89_payload     (clk50Area_keyMatrix_keyStatus_89_payload   ), //o
    .keyStatus_90_valid       (clk50Area_keyMatrix_keyStatus_90_valid     ), //o
    .keyStatus_90_payload     (clk50Area_keyMatrix_keyStatus_90_payload   ), //o
    .keyStatus_91_valid       (clk50Area_keyMatrix_keyStatus_91_valid     ), //o
    .keyStatus_91_payload     (clk50Area_keyMatrix_keyStatus_91_payload   ), //o
    .keyStatus_92_valid       (clk50Area_keyMatrix_keyStatus_92_valid     ), //o
    .keyStatus_92_payload     (clk50Area_keyMatrix_keyStatus_92_payload   ), //o
    .keyStatus_93_valid       (clk50Area_keyMatrix_keyStatus_93_valid     ), //o
    .keyStatus_93_payload     (clk50Area_keyMatrix_keyStatus_93_payload   ), //o
    .keyStatus_94_valid       (clk50Area_keyMatrix_keyStatus_94_valid     ), //o
    .keyStatus_94_payload     (clk50Area_keyMatrix_keyStatus_94_payload   ), //o
    .keyStatus_95_valid       (clk50Area_keyMatrix_keyStatus_95_valid     ), //o
    .keyStatus_95_payload     (clk50Area_keyMatrix_keyStatus_95_payload   ), //o
    .keyStatus_96_valid       (clk50Area_keyMatrix_keyStatus_96_valid     ), //o
    .keyStatus_96_payload     (clk50Area_keyMatrix_keyStatus_96_payload   ), //o
    .keyStatus_97_valid       (clk50Area_keyMatrix_keyStatus_97_valid     ), //o
    .keyStatus_97_payload     (clk50Area_keyMatrix_keyStatus_97_payload   ), //o
    .keyStatus_98_valid       (clk50Area_keyMatrix_keyStatus_98_valid     ), //o
    .keyStatus_98_payload     (clk50Area_keyMatrix_keyStatus_98_payload   ), //o
    .keyStatus_99_valid       (clk50Area_keyMatrix_keyStatus_99_valid     ), //o
    .keyStatus_99_payload     (clk50Area_keyMatrix_keyStatus_99_payload   ), //o
    .keyStatus_100_valid      (clk50Area_keyMatrix_keyStatus_100_valid    ), //o
    .keyStatus_100_payload    (clk50Area_keyMatrix_keyStatus_100_payload  ), //o
    .keyStatus_101_valid      (clk50Area_keyMatrix_keyStatus_101_valid    ), //o
    .keyStatus_101_payload    (clk50Area_keyMatrix_keyStatus_101_payload  ), //o
    .keyStatus_102_valid      (clk50Area_keyMatrix_keyStatus_102_valid    ), //o
    .keyStatus_102_payload    (clk50Area_keyMatrix_keyStatus_102_payload  ), //o
    ._zz_1                    (_zz_1                                      ), //i
    .CLK_50                   (CLK_50                                     )  //i
  );
  UartCtrl uartCtrl_2 (
    .io_config_frame_dataLength    (_zz_8[2:0]                                            ), //i
    .io_config_frame_stop          (_zz_9                                                 ), //i
    .io_config_frame_parity        (_zz_10[1:0]                                           ), //i
    .io_config_clockDivider        (_zz_11[19:0]                                          ), //i
    .io_write_valid                (_zz_3                                                 ), //i
    .io_write_ready                (uartCtrl_2_io_write_ready                             ), //o
    .io_write_payload              (clk50Area_keyMatrix_scanIdx_payload_regNextWhen[7:0]  ), //i
    .io_read_valid                 (uartCtrl_2_io_read_valid                              ), //o
    .io_read_ready                 (_zz_12                                                ), //i
    .io_read_payload               (uartCtrl_2_io_read_payload[7:0]                       ), //o
    .io_uart_txd                   (uartCtrl_2_io_uart_txd                                ), //o
    .io_uart_rxd                   (_zz_13                                                ), //i
    .io_readError                  (uartCtrl_2_io_readError                               ), //o
    .io_writeBreak                 (_zz_14                                                ), //i
    .io_readBreak                  (uartCtrl_2_io_readBreak                               ), //o
    .CLK_50                        (CLK_50                                                ), //i
    ._zz_1                         (_zz_1                                                 )  //i
  );
  HID clk50Area_hid (
    .TXD                      (clk50Area_hid_TXD                         ), //o
    .scanIdx_valid            (clk50Area_keyMatrix_scanIdx_valid         ), //i
    .scanIdx_payload          (clk50Area_keyMatrix_scanIdx_payload[7:0]  ), //i
    .keyStatus_0_valid        (_zz_15                                    ), //i
    .keyStatus_0_payload      (_zz_16                                    ), //i
    .keyStatus_1_valid        (_zz_17                                    ), //i
    .keyStatus_1_payload      (_zz_18                                    ), //i
    .keyStatus_2_valid        (_zz_19                                    ), //i
    .keyStatus_2_payload      (_zz_20                                    ), //i
    .keyStatus_3_valid        (_zz_21                                    ), //i
    .keyStatus_3_payload      (_zz_22                                    ), //i
    .keyStatus_4_valid        (_zz_23                                    ), //i
    .keyStatus_4_payload      (_zz_24                                    ), //i
    .keyStatus_5_valid        (_zz_25                                    ), //i
    .keyStatus_5_payload      (_zz_26                                    ), //i
    .keyStatus_6_valid        (_zz_27                                    ), //i
    .keyStatus_6_payload      (_zz_28                                    ), //i
    .keyStatus_7_valid        (_zz_29                                    ), //i
    .keyStatus_7_payload      (_zz_30                                    ), //i
    .keyStatus_8_valid        (_zz_31                                    ), //i
    .keyStatus_8_payload      (_zz_32                                    ), //i
    .keyStatus_9_valid        (_zz_33                                    ), //i
    .keyStatus_9_payload      (_zz_34                                    ), //i
    .keyStatus_10_valid       (_zz_35                                    ), //i
    .keyStatus_10_payload     (_zz_36                                    ), //i
    .keyStatus_11_valid       (_zz_37                                    ), //i
    .keyStatus_11_payload     (_zz_38                                    ), //i
    .keyStatus_12_valid       (_zz_39                                    ), //i
    .keyStatus_12_payload     (_zz_40                                    ), //i
    .keyStatus_13_valid       (_zz_41                                    ), //i
    .keyStatus_13_payload     (_zz_42                                    ), //i
    .keyStatus_14_valid       (_zz_43                                    ), //i
    .keyStatus_14_payload     (_zz_44                                    ), //i
    .keyStatus_15_valid       (_zz_45                                    ), //i
    .keyStatus_15_payload     (_zz_46                                    ), //i
    .keyStatus_16_valid       (_zz_47                                    ), //i
    .keyStatus_16_payload     (_zz_48                                    ), //i
    .keyStatus_17_valid       (_zz_49                                    ), //i
    .keyStatus_17_payload     (_zz_50                                    ), //i
    .keyStatus_18_valid       (_zz_51                                    ), //i
    .keyStatus_18_payload     (_zz_52                                    ), //i
    .keyStatus_19_valid       (_zz_53                                    ), //i
    .keyStatus_19_payload     (_zz_54                                    ), //i
    .keyStatus_20_valid       (_zz_55                                    ), //i
    .keyStatus_20_payload     (_zz_56                                    ), //i
    .keyStatus_21_valid       (_zz_57                                    ), //i
    .keyStatus_21_payload     (_zz_58                                    ), //i
    .keyStatus_22_valid       (_zz_59                                    ), //i
    .keyStatus_22_payload     (_zz_60                                    ), //i
    .keyStatus_23_valid       (_zz_61                                    ), //i
    .keyStatus_23_payload     (_zz_62                                    ), //i
    .keyStatus_24_valid       (_zz_63                                    ), //i
    .keyStatus_24_payload     (_zz_64                                    ), //i
    .keyStatus_25_valid       (_zz_65                                    ), //i
    .keyStatus_25_payload     (_zz_66                                    ), //i
    .keyStatus_26_valid       (_zz_67                                    ), //i
    .keyStatus_26_payload     (_zz_68                                    ), //i
    .keyStatus_27_valid       (_zz_69                                    ), //i
    .keyStatus_27_payload     (_zz_70                                    ), //i
    .keyStatus_28_valid       (_zz_71                                    ), //i
    .keyStatus_28_payload     (_zz_72                                    ), //i
    .keyStatus_29_valid       (_zz_73                                    ), //i
    .keyStatus_29_payload     (_zz_74                                    ), //i
    .keyStatus_30_valid       (_zz_75                                    ), //i
    .keyStatus_30_payload     (_zz_76                                    ), //i
    .keyStatus_31_valid       (_zz_77                                    ), //i
    .keyStatus_31_payload     (_zz_78                                    ), //i
    .keyStatus_32_valid       (_zz_79                                    ), //i
    .keyStatus_32_payload     (_zz_80                                    ), //i
    .keyStatus_33_valid       (_zz_81                                    ), //i
    .keyStatus_33_payload     (_zz_82                                    ), //i
    .keyStatus_34_valid       (_zz_83                                    ), //i
    .keyStatus_34_payload     (_zz_84                                    ), //i
    .keyStatus_35_valid       (_zz_85                                    ), //i
    .keyStatus_35_payload     (_zz_86                                    ), //i
    .keyStatus_36_valid       (_zz_87                                    ), //i
    .keyStatus_36_payload     (_zz_88                                    ), //i
    .keyStatus_37_valid       (_zz_89                                    ), //i
    .keyStatus_37_payload     (_zz_90                                    ), //i
    .keyStatus_38_valid       (_zz_91                                    ), //i
    .keyStatus_38_payload     (_zz_92                                    ), //i
    .keyStatus_39_valid       (_zz_93                                    ), //i
    .keyStatus_39_payload     (_zz_94                                    ), //i
    .keyStatus_40_valid       (_zz_95                                    ), //i
    .keyStatus_40_payload     (_zz_96                                    ), //i
    .keyStatus_41_valid       (_zz_97                                    ), //i
    .keyStatus_41_payload     (_zz_98                                    ), //i
    .keyStatus_42_valid       (_zz_99                                    ), //i
    .keyStatus_42_payload     (_zz_100                                   ), //i
    .keyStatus_43_valid       (_zz_101                                   ), //i
    .keyStatus_43_payload     (_zz_102                                   ), //i
    .keyStatus_44_valid       (_zz_103                                   ), //i
    .keyStatus_44_payload     (_zz_104                                   ), //i
    .keyStatus_45_valid       (_zz_105                                   ), //i
    .keyStatus_45_payload     (_zz_106                                   ), //i
    .keyStatus_46_valid       (_zz_107                                   ), //i
    .keyStatus_46_payload     (_zz_108                                   ), //i
    .keyStatus_47_valid       (_zz_109                                   ), //i
    .keyStatus_47_payload     (_zz_110                                   ), //i
    .keyStatus_48_valid       (_zz_111                                   ), //i
    .keyStatus_48_payload     (_zz_112                                   ), //i
    .keyStatus_49_valid       (_zz_113                                   ), //i
    .keyStatus_49_payload     (_zz_114                                   ), //i
    .keyStatus_50_valid       (_zz_115                                   ), //i
    .keyStatus_50_payload     (_zz_116                                   ), //i
    .keyStatus_51_valid       (_zz_117                                   ), //i
    .keyStatus_51_payload     (_zz_118                                   ), //i
    .keyStatus_52_valid       (_zz_119                                   ), //i
    .keyStatus_52_payload     (_zz_120                                   ), //i
    .keyStatus_53_valid       (_zz_121                                   ), //i
    .keyStatus_53_payload     (_zz_122                                   ), //i
    .keyStatus_54_valid       (_zz_123                                   ), //i
    .keyStatus_54_payload     (_zz_124                                   ), //i
    .keyStatus_55_valid       (_zz_125                                   ), //i
    .keyStatus_55_payload     (_zz_126                                   ), //i
    .keyStatus_56_valid       (_zz_127                                   ), //i
    .keyStatus_56_payload     (_zz_128                                   ), //i
    .keyStatus_57_valid       (_zz_129                                   ), //i
    .keyStatus_57_payload     (_zz_130                                   ), //i
    .keyStatus_58_valid       (_zz_131                                   ), //i
    .keyStatus_58_payload     (_zz_132                                   ), //i
    .keyStatus_59_valid       (_zz_133                                   ), //i
    .keyStatus_59_payload     (_zz_134                                   ), //i
    .keyStatus_60_valid       (_zz_135                                   ), //i
    .keyStatus_60_payload     (_zz_136                                   ), //i
    .keyStatus_61_valid       (_zz_137                                   ), //i
    .keyStatus_61_payload     (_zz_138                                   ), //i
    .keyStatus_62_valid       (_zz_139                                   ), //i
    .keyStatus_62_payload     (_zz_140                                   ), //i
    .keyStatus_63_valid       (_zz_141                                   ), //i
    .keyStatus_63_payload     (_zz_142                                   ), //i
    .keyStatus_64_valid       (_zz_143                                   ), //i
    .keyStatus_64_payload     (_zz_144                                   ), //i
    .keyStatus_65_valid       (_zz_145                                   ), //i
    .keyStatus_65_payload     (_zz_146                                   ), //i
    .keyStatus_66_valid       (_zz_147                                   ), //i
    .keyStatus_66_payload     (_zz_148                                   ), //i
    .keyStatus_67_valid       (_zz_149                                   ), //i
    .keyStatus_67_payload     (_zz_150                                   ), //i
    .keyStatus_68_valid       (_zz_151                                   ), //i
    .keyStatus_68_payload     (_zz_152                                   ), //i
    .keyStatus_69_valid       (_zz_153                                   ), //i
    .keyStatus_69_payload     (_zz_154                                   ), //i
    .keyStatus_70_valid       (_zz_155                                   ), //i
    .keyStatus_70_payload     (_zz_156                                   ), //i
    .keyStatus_71_valid       (_zz_157                                   ), //i
    .keyStatus_71_payload     (_zz_158                                   ), //i
    .keyStatus_72_valid       (_zz_159                                   ), //i
    .keyStatus_72_payload     (_zz_160                                   ), //i
    .keyStatus_73_valid       (_zz_161                                   ), //i
    .keyStatus_73_payload     (_zz_162                                   ), //i
    .keyStatus_74_valid       (clk50Area_keyMatrix_keyStatus_74_valid    ), //i
    .keyStatus_74_payload     (clk50Area_keyMatrix_keyStatus_74_payload  ), //i
    .keyStatus_75_valid       (_zz_163                                   ), //i
    .keyStatus_75_payload     (_zz_164                                   ), //i
    .keyStatus_76_valid       (_zz_165                                   ), //i
    .keyStatus_76_payload     (_zz_166                                   ), //i
    .keyStatus_77_valid       (_zz_167                                   ), //i
    .keyStatus_77_payload     (_zz_168                                   ), //i
    .keyStatus_78_valid       (_zz_169                                   ), //i
    .keyStatus_78_payload     (_zz_170                                   ), //i
    .keyStatus_79_valid       (_zz_171                                   ), //i
    .keyStatus_79_payload     (_zz_172                                   ), //i
    .keyStatus_80_valid       (_zz_173                                   ), //i
    .keyStatus_80_payload     (_zz_174                                   ), //i
    .keyStatus_81_valid       (_zz_175                                   ), //i
    .keyStatus_81_payload     (_zz_176                                   ), //i
    .keyStatus_82_valid       (_zz_177                                   ), //i
    .keyStatus_82_payload     (_zz_178                                   ), //i
    .keyStatus_83_valid       (_zz_179                                   ), //i
    .keyStatus_83_payload     (_zz_180                                   ), //i
    .keyStatus_84_valid       (_zz_181                                   ), //i
    .keyStatus_84_payload     (_zz_182                                   ), //i
    .keyStatus_85_valid       (clk50Area_keyMatrix_keyStatus_85_valid    ), //i
    .keyStatus_85_payload     (clk50Area_keyMatrix_keyStatus_85_payload  ), //i
    .keyStatus_86_valid       (_zz_183                                   ), //i
    .keyStatus_86_payload     (_zz_184                                   ), //i
    .keyStatus_87_valid       (_zz_185                                   ), //i
    .keyStatus_87_payload     (_zz_186                                   ), //i
    .keyStatus_88_valid       (_zz_187                                   ), //i
    .keyStatus_88_payload     (_zz_188                                   ), //i
    .keyStatus_89_valid       (_zz_189                                   ), //i
    .keyStatus_89_payload     (_zz_190                                   ), //i
    .keyStatus_90_valid       (clk50Area_keyMatrix_keyStatus_90_valid    ), //i
    .keyStatus_90_payload     (clk50Area_keyMatrix_keyStatus_90_payload  ), //i
    .keyStatus_91_valid       (clk50Area_keyMatrix_keyStatus_91_valid    ), //i
    .keyStatus_91_payload     (clk50Area_keyMatrix_keyStatus_91_payload  ), //i
    .keyStatus_92_valid       (clk50Area_keyMatrix_keyStatus_92_valid    ), //i
    .keyStatus_92_payload     (clk50Area_keyMatrix_keyStatus_92_payload  ), //i
    .keyStatus_93_valid       (_zz_191                                   ), //i
    .keyStatus_93_payload     (_zz_192                                   ), //i
    .keyStatus_94_valid       (clk50Area_keyMatrix_keyStatus_94_valid    ), //i
    .keyStatus_94_payload     (clk50Area_keyMatrix_keyStatus_94_payload  ), //i
    .keyStatus_95_valid       (_zz_193                                   ), //i
    .keyStatus_95_payload     (_zz_194                                   ), //i
    .keyStatus_96_valid       (clk50Area_keyMatrix_keyStatus_96_valid    ), //i
    .keyStatus_96_payload     (clk50Area_keyMatrix_keyStatus_96_payload  ), //i
    .keyStatus_97_valid       (_zz_195                                   ), //i
    .keyStatus_97_payload     (_zz_196                                   ), //i
    .keyStatus_98_valid       (_zz_197                                   ), //i
    .keyStatus_98_payload     (_zz_198                                   ), //i
    .keyStatus_99_valid       (_zz_199                                   ), //i
    .keyStatus_99_payload     (_zz_200                                   ), //i
    .keyStatus_100_valid      (_zz_201                                   ), //i
    .keyStatus_100_payload    (_zz_202                                   ), //i
    .keyStatus_101_valid      (_zz_203                                   ), //i
    .keyStatus_101_payload    (_zz_204                                   ), //i
    .keyStatus_102_valid      (_zz_205                                   ), //i
    .keyStatus_102_payload    (_zz_206                                   ), //i
    .CLK_50                   (CLK_50                                    ), //i
    ._zz_1                    (_zz_1                                     )  //i
  );
  assign _zz_4 = (! KEY_Fn);
  always @ (*) begin
    _zz_1 = 1'b0;
    _zz_1 = bufferCC_3_io_dataOut;
  end

  assign _zz_2 = (rstCtrl_io_globalReset || (! pll100_locked));
  assign _zz_5 = 1'b0;
  assign _zz_6 = (! _zz_1);
  assign LED_A = core_io_row;
  assign LED_K = core_io_col;
  assign flash_dclk = core_flash_dclk;
  assign flash_sce = core_flash_sce;
  assign flash_sdo = core_flash_sdo;
  assign LED_R6 = _zz_1;
  assign ROW = clk50Area_keyMatrix_ROW;
  assign _zz_7 = 1'b1;
  assign _zz_11 = 20'h00035;
  assign _zz_8 = 3'b111;
  assign _zz_10 = `UartParityType_defaultEncoding_NONE;
  assign _zz_9 = `UartStopType_defaultEncoding_ONE;
  assign _zz_14 = 1'b0;
  assign _zz_13 = 1'b1;
  assign TXD = clk50Area_hid_TXD;
  always @ (posedge CLK_50) begin
    if(clk50Area_keyMatrix_scanIdx_valid)begin
      clk50Area_keyMatrix_scanIdx_payload_regNextWhen <= clk50Area_keyMatrix_scanIdx_payload;
    end
  end

  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      _zz_3 <= 1'b0;
    end else begin
      if(clk50Area_keyMatrix_scanIdx_valid)begin
        _zz_3 <= 1'b1;
      end else begin
        if(uartCtrl_2_io_write_ready)begin
          _zz_3 <= 1'b0;
        end
      end
    end
  end


endmodule

module HID (
  output              TXD,
  input               scanIdx_valid,
  input      [7:0]    scanIdx_payload,
  input               keyStatus_0_valid,
  input               keyStatus_0_payload,
  input               keyStatus_1_valid,
  input               keyStatus_1_payload,
  input               keyStatus_2_valid,
  input               keyStatus_2_payload,
  input               keyStatus_3_valid,
  input               keyStatus_3_payload,
  input               keyStatus_4_valid,
  input               keyStatus_4_payload,
  input               keyStatus_5_valid,
  input               keyStatus_5_payload,
  input               keyStatus_6_valid,
  input               keyStatus_6_payload,
  input               keyStatus_7_valid,
  input               keyStatus_7_payload,
  input               keyStatus_8_valid,
  input               keyStatus_8_payload,
  input               keyStatus_9_valid,
  input               keyStatus_9_payload,
  input               keyStatus_10_valid,
  input               keyStatus_10_payload,
  input               keyStatus_11_valid,
  input               keyStatus_11_payload,
  input               keyStatus_12_valid,
  input               keyStatus_12_payload,
  input               keyStatus_13_valid,
  input               keyStatus_13_payload,
  input               keyStatus_14_valid,
  input               keyStatus_14_payload,
  input               keyStatus_15_valid,
  input               keyStatus_15_payload,
  input               keyStatus_16_valid,
  input               keyStatus_16_payload,
  input               keyStatus_17_valid,
  input               keyStatus_17_payload,
  input               keyStatus_18_valid,
  input               keyStatus_18_payload,
  input               keyStatus_19_valid,
  input               keyStatus_19_payload,
  input               keyStatus_20_valid,
  input               keyStatus_20_payload,
  input               keyStatus_21_valid,
  input               keyStatus_21_payload,
  input               keyStatus_22_valid,
  input               keyStatus_22_payload,
  input               keyStatus_23_valid,
  input               keyStatus_23_payload,
  input               keyStatus_24_valid,
  input               keyStatus_24_payload,
  input               keyStatus_25_valid,
  input               keyStatus_25_payload,
  input               keyStatus_26_valid,
  input               keyStatus_26_payload,
  input               keyStatus_27_valid,
  input               keyStatus_27_payload,
  input               keyStatus_28_valid,
  input               keyStatus_28_payload,
  input               keyStatus_29_valid,
  input               keyStatus_29_payload,
  input               keyStatus_30_valid,
  input               keyStatus_30_payload,
  input               keyStatus_31_valid,
  input               keyStatus_31_payload,
  input               keyStatus_32_valid,
  input               keyStatus_32_payload,
  input               keyStatus_33_valid,
  input               keyStatus_33_payload,
  input               keyStatus_34_valid,
  input               keyStatus_34_payload,
  input               keyStatus_35_valid,
  input               keyStatus_35_payload,
  input               keyStatus_36_valid,
  input               keyStatus_36_payload,
  input               keyStatus_37_valid,
  input               keyStatus_37_payload,
  input               keyStatus_38_valid,
  input               keyStatus_38_payload,
  input               keyStatus_39_valid,
  input               keyStatus_39_payload,
  input               keyStatus_40_valid,
  input               keyStatus_40_payload,
  input               keyStatus_41_valid,
  input               keyStatus_41_payload,
  input               keyStatus_42_valid,
  input               keyStatus_42_payload,
  input               keyStatus_43_valid,
  input               keyStatus_43_payload,
  input               keyStatus_44_valid,
  input               keyStatus_44_payload,
  input               keyStatus_45_valid,
  input               keyStatus_45_payload,
  input               keyStatus_46_valid,
  input               keyStatus_46_payload,
  input               keyStatus_47_valid,
  input               keyStatus_47_payload,
  input               keyStatus_48_valid,
  input               keyStatus_48_payload,
  input               keyStatus_49_valid,
  input               keyStatus_49_payload,
  input               keyStatus_50_valid,
  input               keyStatus_50_payload,
  input               keyStatus_51_valid,
  input               keyStatus_51_payload,
  input               keyStatus_52_valid,
  input               keyStatus_52_payload,
  input               keyStatus_53_valid,
  input               keyStatus_53_payload,
  input               keyStatus_54_valid,
  input               keyStatus_54_payload,
  input               keyStatus_55_valid,
  input               keyStatus_55_payload,
  input               keyStatus_56_valid,
  input               keyStatus_56_payload,
  input               keyStatus_57_valid,
  input               keyStatus_57_payload,
  input               keyStatus_58_valid,
  input               keyStatus_58_payload,
  input               keyStatus_59_valid,
  input               keyStatus_59_payload,
  input               keyStatus_60_valid,
  input               keyStatus_60_payload,
  input               keyStatus_61_valid,
  input               keyStatus_61_payload,
  input               keyStatus_62_valid,
  input               keyStatus_62_payload,
  input               keyStatus_63_valid,
  input               keyStatus_63_payload,
  input               keyStatus_64_valid,
  input               keyStatus_64_payload,
  input               keyStatus_65_valid,
  input               keyStatus_65_payload,
  input               keyStatus_66_valid,
  input               keyStatus_66_payload,
  input               keyStatus_67_valid,
  input               keyStatus_67_payload,
  input               keyStatus_68_valid,
  input               keyStatus_68_payload,
  input               keyStatus_69_valid,
  input               keyStatus_69_payload,
  input               keyStatus_70_valid,
  input               keyStatus_70_payload,
  input               keyStatus_71_valid,
  input               keyStatus_71_payload,
  input               keyStatus_72_valid,
  input               keyStatus_72_payload,
  input               keyStatus_73_valid,
  input               keyStatus_73_payload,
  input               keyStatus_74_valid,
  input               keyStatus_74_payload,
  input               keyStatus_75_valid,
  input               keyStatus_75_payload,
  input               keyStatus_76_valid,
  input               keyStatus_76_payload,
  input               keyStatus_77_valid,
  input               keyStatus_77_payload,
  input               keyStatus_78_valid,
  input               keyStatus_78_payload,
  input               keyStatus_79_valid,
  input               keyStatus_79_payload,
  input               keyStatus_80_valid,
  input               keyStatus_80_payload,
  input               keyStatus_81_valid,
  input               keyStatus_81_payload,
  input               keyStatus_82_valid,
  input               keyStatus_82_payload,
  input               keyStatus_83_valid,
  input               keyStatus_83_payload,
  input               keyStatus_84_valid,
  input               keyStatus_84_payload,
  input               keyStatus_85_valid,
  input               keyStatus_85_payload,
  input               keyStatus_86_valid,
  input               keyStatus_86_payload,
  input               keyStatus_87_valid,
  input               keyStatus_87_payload,
  input               keyStatus_88_valid,
  input               keyStatus_88_payload,
  input               keyStatus_89_valid,
  input               keyStatus_89_payload,
  input               keyStatus_90_valid,
  input               keyStatus_90_payload,
  input               keyStatus_91_valid,
  input               keyStatus_91_payload,
  input               keyStatus_92_valid,
  input               keyStatus_92_payload,
  input               keyStatus_93_valid,
  input               keyStatus_93_payload,
  input               keyStatus_94_valid,
  input               keyStatus_94_payload,
  input               keyStatus_95_valid,
  input               keyStatus_95_payload,
  input               keyStatus_96_valid,
  input               keyStatus_96_payload,
  input               keyStatus_97_valid,
  input               keyStatus_97_payload,
  input               keyStatus_98_valid,
  input               keyStatus_98_payload,
  input               keyStatus_99_valid,
  input               keyStatus_99_payload,
  input               keyStatus_100_valid,
  input               keyStatus_100_payload,
  input               keyStatus_101_valid,
  input               keyStatus_101_payload,
  input               keyStatus_102_valid,
  input               keyStatus_102_payload,
  input               CLK_50,
  input               _zz_1
);
  wire       [2:0]    _zz_2;
  wire       `UartStopType_defaultEncoding_type _zz_3;
  wire       `UartParityType_defaultEncoding_type _zz_4;
  wire       [19:0]   _zz_5;
  wire                _zz_6;
  reg        [7:0]    _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  reg        [7:0]    _zz_11;
  wire                uartCtrl_2_io_write_ready;
  wire                uartCtrl_2_io_read_valid;
  wire       [7:0]    uartCtrl_2_io_read_payload;
  wire                uartCtrl_2_io_uart_txd;
  wire                uartCtrl_2_io_readError;
  wire                uartCtrl_2_io_readBreak;
  wire                _zz_12;
  reg        [6:0]    idxLatch;
  reg                 staLatch;
  wire                machine_wantExit;
  reg                 machine_wantStart;
  reg        `machine_enumDefinition_defaultEncoding_type machine_stateReg;
  reg        `machine_enumDefinition_defaultEncoding_type machine_stateNext;
  `ifndef SYNTHESIS
  reg [127:0] machine_stateReg_string;
  reg [127:0] machine_stateNext_string;
  `endif

  (* ram_init_file = "VerilogHDL/hid.mif" *) reg [7:0] hidKeyTable [0:127];

  assign _zz_12 = 1'b1;
  always @ (posedge CLK_50) begin
    if(_zz_12) begin
      _zz_11 <= hidKeyTable[idxLatch];
    end
  end

  UartCtrl uartCtrl_2 (
    .io_config_frame_dataLength    (_zz_2[2:0]                       ), //i
    .io_config_frame_stop          (_zz_3                            ), //i
    .io_config_frame_parity        (_zz_4[1:0]                       ), //i
    .io_config_clockDivider        (_zz_5[19:0]                      ), //i
    .io_write_valid                (_zz_6                            ), //i
    .io_write_ready                (uartCtrl_2_io_write_ready        ), //o
    .io_write_payload              (_zz_7[7:0]                       ), //i
    .io_read_valid                 (uartCtrl_2_io_read_valid         ), //o
    .io_read_ready                 (_zz_8                            ), //i
    .io_read_payload               (uartCtrl_2_io_read_payload[7:0]  ), //o
    .io_uart_txd                   (uartCtrl_2_io_uart_txd           ), //o
    .io_uart_rxd                   (_zz_9                            ), //i
    .io_readError                  (uartCtrl_2_io_readError          ), //o
    .io_writeBreak                 (_zz_10                           ), //i
    .io_readBreak                  (uartCtrl_2_io_readBreak          ), //o
    .CLK_50                        (CLK_50                           ), //i
    ._zz_1                         (_zz_1                            )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_BOOT : machine_stateReg_string = "machine_BOOT    ";
      `machine_enumDefinition_defaultEncoding_machine_idle : machine_stateReg_string = "machine_idle    ";
      `machine_enumDefinition_defaultEncoding_machine_k6 : machine_stateReg_string = "machine_k6      ";
      `machine_enumDefinition_defaultEncoding_machine_k5 : machine_stateReg_string = "machine_k5      ";
      `machine_enumDefinition_defaultEncoding_machine_k4 : machine_stateReg_string = "machine_k4      ";
      `machine_enumDefinition_defaultEncoding_machine_k3 : machine_stateReg_string = "machine_k3      ";
      `machine_enumDefinition_defaultEncoding_machine_k2 : machine_stateReg_string = "machine_k2      ";
      `machine_enumDefinition_defaultEncoding_machine_k1 : machine_stateReg_string = "machine_k1      ";
      `machine_enumDefinition_defaultEncoding_machine_reserved : machine_stateReg_string = "machine_reserved";
      `machine_enumDefinition_defaultEncoding_machine_special : machine_stateReg_string = "machine_special ";
      default : machine_stateReg_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(machine_stateNext)
      `machine_enumDefinition_defaultEncoding_machine_BOOT : machine_stateNext_string = "machine_BOOT    ";
      `machine_enumDefinition_defaultEncoding_machine_idle : machine_stateNext_string = "machine_idle    ";
      `machine_enumDefinition_defaultEncoding_machine_k6 : machine_stateNext_string = "machine_k6      ";
      `machine_enumDefinition_defaultEncoding_machine_k5 : machine_stateNext_string = "machine_k5      ";
      `machine_enumDefinition_defaultEncoding_machine_k4 : machine_stateNext_string = "machine_k4      ";
      `machine_enumDefinition_defaultEncoding_machine_k3 : machine_stateNext_string = "machine_k3      ";
      `machine_enumDefinition_defaultEncoding_machine_k2 : machine_stateNext_string = "machine_k2      ";
      `machine_enumDefinition_defaultEncoding_machine_k1 : machine_stateNext_string = "machine_k1      ";
      `machine_enumDefinition_defaultEncoding_machine_reserved : machine_stateNext_string = "machine_reserved";
      `machine_enumDefinition_defaultEncoding_machine_special : machine_stateNext_string = "machine_special ";
      default : machine_stateNext_string = "????????????????";
    endcase
  end
  `endif

  assign _zz_5 = 20'h0028a;
  assign _zz_2 = 3'b111;
  assign _zz_4 = `UartParityType_defaultEncoding_NONE;
  assign _zz_3 = `UartStopType_defaultEncoding_ONE;
  assign _zz_9 = 1'b1;
  assign _zz_10 = 1'b0;
  always @ (*) begin
    _zz_7 = 8'h0;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k6 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k5 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k4 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k3 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k2 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k1 : begin
        if(staLatch)begin
          _zz_7 = _zz_11;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_reserved : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_special : begin
        _zz_7 = {1'b0,{keyStatus_94_payload,{keyStatus_85_payload,{keyStatus_96_payload,{keyStatus_91_payload,{keyStatus_92_payload,{keyStatus_74_payload,keyStatus_90_payload}}}}}}};
      end
      default : begin
      end
    endcase
  end

  assign TXD = uartCtrl_2_io_uart_txd;
  assign machine_wantExit = 1'b0;
  always @ (*) begin
    machine_wantStart = 1'b0;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k6 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k5 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k4 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k3 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k2 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_k1 : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_reserved : begin
      end
      `machine_enumDefinition_defaultEncoding_machine_special : begin
      end
      default : begin
        machine_wantStart = 1'b1;
      end
    endcase
  end

  assign _zz_6 = (! (machine_stateReg == `machine_enumDefinition_defaultEncoding_machine_idle));
  always @ (*) begin
    machine_stateNext = machine_stateReg;
    case(machine_stateReg)
      `machine_enumDefinition_defaultEncoding_machine_idle : begin
        if(scanIdx_valid)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_special;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_k6 : begin
        if(uartCtrl_2_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_idle;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_k5 : begin
        if(uartCtrl_2_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_k6;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_k4 : begin
        if(uartCtrl_2_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_k5;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_k3 : begin
        if(uartCtrl_2_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_k4;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_k2 : begin
        if(uartCtrl_2_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_k3;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_k1 : begin
        if(uartCtrl_2_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_k2;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_reserved : begin
        if(uartCtrl_2_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_k1;
        end
      end
      `machine_enumDefinition_defaultEncoding_machine_special : begin
        if(uartCtrl_2_io_write_ready)begin
          machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_reserved;
        end
      end
      default : begin
      end
    endcase
    if(machine_wantStart)begin
      machine_stateNext = `machine_enumDefinition_defaultEncoding_machine_idle;
    end
  end

  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      idxLatch <= 7'h0;
      staLatch <= 1'b0;
      machine_stateReg <= `machine_enumDefinition_defaultEncoding_machine_BOOT;
    end else begin
      if(scanIdx_valid)begin
        idxLatch <= scanIdx_payload[6 : 0];
      end
      if(scanIdx_valid)begin
        staLatch <= scanIdx_payload[7];
      end
      machine_stateReg <= machine_stateNext;
    end
  end


endmodule

//UartCtrl replaced by UartCtrl

module KeyMatrix (
  input               enabled,
  input      [20:0]   COL,
  output     [5:0]    ROW,
  output              scanIdx_valid,
  output     [7:0]    scanIdx_payload,
  output              keyStatus_0_valid,
  output              keyStatus_0_payload,
  output              keyStatus_1_valid,
  output              keyStatus_1_payload,
  output              keyStatus_2_valid,
  output              keyStatus_2_payload,
  output              keyStatus_3_valid,
  output              keyStatus_3_payload,
  output              keyStatus_4_valid,
  output              keyStatus_4_payload,
  output              keyStatus_5_valid,
  output              keyStatus_5_payload,
  output              keyStatus_6_valid,
  output              keyStatus_6_payload,
  output              keyStatus_7_valid,
  output              keyStatus_7_payload,
  output              keyStatus_8_valid,
  output              keyStatus_8_payload,
  output              keyStatus_9_valid,
  output              keyStatus_9_payload,
  output              keyStatus_10_valid,
  output              keyStatus_10_payload,
  output              keyStatus_11_valid,
  output              keyStatus_11_payload,
  output              keyStatus_12_valid,
  output              keyStatus_12_payload,
  output              keyStatus_13_valid,
  output              keyStatus_13_payload,
  output              keyStatus_14_valid,
  output              keyStatus_14_payload,
  output              keyStatus_15_valid,
  output              keyStatus_15_payload,
  output              keyStatus_16_valid,
  output              keyStatus_16_payload,
  output              keyStatus_17_valid,
  output              keyStatus_17_payload,
  output              keyStatus_18_valid,
  output              keyStatus_18_payload,
  output              keyStatus_19_valid,
  output              keyStatus_19_payload,
  output              keyStatus_20_valid,
  output              keyStatus_20_payload,
  output              keyStatus_21_valid,
  output              keyStatus_21_payload,
  output              keyStatus_22_valid,
  output              keyStatus_22_payload,
  output              keyStatus_23_valid,
  output              keyStatus_23_payload,
  output              keyStatus_24_valid,
  output              keyStatus_24_payload,
  output              keyStatus_25_valid,
  output              keyStatus_25_payload,
  output              keyStatus_26_valid,
  output              keyStatus_26_payload,
  output              keyStatus_27_valid,
  output              keyStatus_27_payload,
  output              keyStatus_28_valid,
  output              keyStatus_28_payload,
  output              keyStatus_29_valid,
  output              keyStatus_29_payload,
  output              keyStatus_30_valid,
  output              keyStatus_30_payload,
  output              keyStatus_31_valid,
  output              keyStatus_31_payload,
  output              keyStatus_32_valid,
  output              keyStatus_32_payload,
  output              keyStatus_33_valid,
  output              keyStatus_33_payload,
  output              keyStatus_34_valid,
  output              keyStatus_34_payload,
  output              keyStatus_35_valid,
  output              keyStatus_35_payload,
  output              keyStatus_36_valid,
  output              keyStatus_36_payload,
  output              keyStatus_37_valid,
  output              keyStatus_37_payload,
  output              keyStatus_38_valid,
  output              keyStatus_38_payload,
  output              keyStatus_39_valid,
  output              keyStatus_39_payload,
  output              keyStatus_40_valid,
  output              keyStatus_40_payload,
  output              keyStatus_41_valid,
  output              keyStatus_41_payload,
  output              keyStatus_42_valid,
  output              keyStatus_42_payload,
  output              keyStatus_43_valid,
  output              keyStatus_43_payload,
  output              keyStatus_44_valid,
  output              keyStatus_44_payload,
  output              keyStatus_45_valid,
  output              keyStatus_45_payload,
  output              keyStatus_46_valid,
  output              keyStatus_46_payload,
  output              keyStatus_47_valid,
  output              keyStatus_47_payload,
  output              keyStatus_48_valid,
  output              keyStatus_48_payload,
  output              keyStatus_49_valid,
  output              keyStatus_49_payload,
  output              keyStatus_50_valid,
  output              keyStatus_50_payload,
  output              keyStatus_51_valid,
  output              keyStatus_51_payload,
  output              keyStatus_52_valid,
  output              keyStatus_52_payload,
  output              keyStatus_53_valid,
  output              keyStatus_53_payload,
  output              keyStatus_54_valid,
  output              keyStatus_54_payload,
  output              keyStatus_55_valid,
  output              keyStatus_55_payload,
  output              keyStatus_56_valid,
  output              keyStatus_56_payload,
  output              keyStatus_57_valid,
  output              keyStatus_57_payload,
  output              keyStatus_58_valid,
  output              keyStatus_58_payload,
  output              keyStatus_59_valid,
  output              keyStatus_59_payload,
  output              keyStatus_60_valid,
  output              keyStatus_60_payload,
  output              keyStatus_61_valid,
  output              keyStatus_61_payload,
  output              keyStatus_62_valid,
  output              keyStatus_62_payload,
  output              keyStatus_63_valid,
  output              keyStatus_63_payload,
  output              keyStatus_64_valid,
  output              keyStatus_64_payload,
  output              keyStatus_65_valid,
  output              keyStatus_65_payload,
  output              keyStatus_66_valid,
  output              keyStatus_66_payload,
  output              keyStatus_67_valid,
  output              keyStatus_67_payload,
  output              keyStatus_68_valid,
  output              keyStatus_68_payload,
  output              keyStatus_69_valid,
  output              keyStatus_69_payload,
  output              keyStatus_70_valid,
  output              keyStatus_70_payload,
  output              keyStatus_71_valid,
  output              keyStatus_71_payload,
  output              keyStatus_72_valid,
  output              keyStatus_72_payload,
  output              keyStatus_73_valid,
  output              keyStatus_73_payload,
  output              keyStatus_74_valid,
  output              keyStatus_74_payload,
  output              keyStatus_75_valid,
  output              keyStatus_75_payload,
  output              keyStatus_76_valid,
  output              keyStatus_76_payload,
  output              keyStatus_77_valid,
  output              keyStatus_77_payload,
  output              keyStatus_78_valid,
  output              keyStatus_78_payload,
  output              keyStatus_79_valid,
  output              keyStatus_79_payload,
  output              keyStatus_80_valid,
  output              keyStatus_80_payload,
  output              keyStatus_81_valid,
  output              keyStatus_81_payload,
  output              keyStatus_82_valid,
  output              keyStatus_82_payload,
  output              keyStatus_83_valid,
  output              keyStatus_83_payload,
  output              keyStatus_84_valid,
  output              keyStatus_84_payload,
  output              keyStatus_85_valid,
  output              keyStatus_85_payload,
  output              keyStatus_86_valid,
  output              keyStatus_86_payload,
  output              keyStatus_87_valid,
  output              keyStatus_87_payload,
  output              keyStatus_88_valid,
  output              keyStatus_88_payload,
  output              keyStatus_89_valid,
  output              keyStatus_89_payload,
  output              keyStatus_90_valid,
  output              keyStatus_90_payload,
  output              keyStatus_91_valid,
  output              keyStatus_91_payload,
  output              keyStatus_92_valid,
  output              keyStatus_92_payload,
  output              keyStatus_93_valid,
  output              keyStatus_93_payload,
  output              keyStatus_94_valid,
  output              keyStatus_94_payload,
  output              keyStatus_95_valid,
  output              keyStatus_95_payload,
  output              keyStatus_96_valid,
  output              keyStatus_96_payload,
  output              keyStatus_97_valid,
  output              keyStatus_97_payload,
  output              keyStatus_98_valid,
  output              keyStatus_98_payload,
  output              keyStatus_99_valid,
  output              keyStatus_99_payload,
  output              keyStatus_100_valid,
  output              keyStatus_100_payload,
  output              keyStatus_101_valid,
  output              keyStatus_101_payload,
  output              keyStatus_102_valid,
  output              keyStatus_102_payload,
  input               _zz_1,
  input               CLK_50
);
  reg                 _zz_9;
  reg                 _zz_10;
  wire       [5:0]    scanK_ROW;
  wire       [102:0]  scanK_key_down;
  wire                debounce_1_keyStatus_0_valid;
  wire                debounce_1_keyStatus_0_payload;
  wire                debounce_1_keyStatus_1_valid;
  wire                debounce_1_keyStatus_1_payload;
  wire                debounce_1_keyStatus_2_valid;
  wire                debounce_1_keyStatus_2_payload;
  wire                debounce_1_keyStatus_3_valid;
  wire                debounce_1_keyStatus_3_payload;
  wire                debounce_1_keyStatus_4_valid;
  wire                debounce_1_keyStatus_4_payload;
  wire                debounce_1_keyStatus_5_valid;
  wire                debounce_1_keyStatus_5_payload;
  wire                debounce_1_keyStatus_6_valid;
  wire                debounce_1_keyStatus_6_payload;
  wire                debounce_1_keyStatus_7_valid;
  wire                debounce_1_keyStatus_7_payload;
  wire                debounce_1_keyStatus_8_valid;
  wire                debounce_1_keyStatus_8_payload;
  wire                debounce_1_keyStatus_9_valid;
  wire                debounce_1_keyStatus_9_payload;
  wire                debounce_1_keyStatus_10_valid;
  wire                debounce_1_keyStatus_10_payload;
  wire                debounce_1_keyStatus_11_valid;
  wire                debounce_1_keyStatus_11_payload;
  wire                debounce_1_keyStatus_12_valid;
  wire                debounce_1_keyStatus_12_payload;
  wire                debounce_1_keyStatus_13_valid;
  wire                debounce_1_keyStatus_13_payload;
  wire                debounce_1_keyStatus_14_valid;
  wire                debounce_1_keyStatus_14_payload;
  wire                debounce_1_keyStatus_15_valid;
  wire                debounce_1_keyStatus_15_payload;
  wire                debounce_1_keyStatus_16_valid;
  wire                debounce_1_keyStatus_16_payload;
  wire                debounce_1_keyStatus_17_valid;
  wire                debounce_1_keyStatus_17_payload;
  wire                debounce_1_keyStatus_18_valid;
  wire                debounce_1_keyStatus_18_payload;
  wire                debounce_1_keyStatus_19_valid;
  wire                debounce_1_keyStatus_19_payload;
  wire                debounce_1_keyStatus_20_valid;
  wire                debounce_1_keyStatus_20_payload;
  wire                debounce_1_keyStatus_21_valid;
  wire                debounce_1_keyStatus_21_payload;
  wire                debounce_1_keyStatus_22_valid;
  wire                debounce_1_keyStatus_22_payload;
  wire                debounce_1_keyStatus_23_valid;
  wire                debounce_1_keyStatus_23_payload;
  wire                debounce_1_keyStatus_24_valid;
  wire                debounce_1_keyStatus_24_payload;
  wire                debounce_1_keyStatus_25_valid;
  wire                debounce_1_keyStatus_25_payload;
  wire                debounce_1_keyStatus_26_valid;
  wire                debounce_1_keyStatus_26_payload;
  wire                debounce_1_keyStatus_27_valid;
  wire                debounce_1_keyStatus_27_payload;
  wire                debounce_1_keyStatus_28_valid;
  wire                debounce_1_keyStatus_28_payload;
  wire                debounce_1_keyStatus_29_valid;
  wire                debounce_1_keyStatus_29_payload;
  wire                debounce_1_keyStatus_30_valid;
  wire                debounce_1_keyStatus_30_payload;
  wire                debounce_1_keyStatus_31_valid;
  wire                debounce_1_keyStatus_31_payload;
  wire                debounce_1_keyStatus_32_valid;
  wire                debounce_1_keyStatus_32_payload;
  wire                debounce_1_keyStatus_33_valid;
  wire                debounce_1_keyStatus_33_payload;
  wire                debounce_1_keyStatus_34_valid;
  wire                debounce_1_keyStatus_34_payload;
  wire                debounce_1_keyStatus_35_valid;
  wire                debounce_1_keyStatus_35_payload;
  wire                debounce_1_keyStatus_36_valid;
  wire                debounce_1_keyStatus_36_payload;
  wire                debounce_1_keyStatus_37_valid;
  wire                debounce_1_keyStatus_37_payload;
  wire                debounce_1_keyStatus_38_valid;
  wire                debounce_1_keyStatus_38_payload;
  wire                debounce_1_keyStatus_39_valid;
  wire                debounce_1_keyStatus_39_payload;
  wire                debounce_1_keyStatus_40_valid;
  wire                debounce_1_keyStatus_40_payload;
  wire                debounce_1_keyStatus_41_valid;
  wire                debounce_1_keyStatus_41_payload;
  wire                debounce_1_keyStatus_42_valid;
  wire                debounce_1_keyStatus_42_payload;
  wire                debounce_1_keyStatus_43_valid;
  wire                debounce_1_keyStatus_43_payload;
  wire                debounce_1_keyStatus_44_valid;
  wire                debounce_1_keyStatus_44_payload;
  wire                debounce_1_keyStatus_45_valid;
  wire                debounce_1_keyStatus_45_payload;
  wire                debounce_1_keyStatus_46_valid;
  wire                debounce_1_keyStatus_46_payload;
  wire                debounce_1_keyStatus_47_valid;
  wire                debounce_1_keyStatus_47_payload;
  wire                debounce_1_keyStatus_48_valid;
  wire                debounce_1_keyStatus_48_payload;
  wire                debounce_1_keyStatus_49_valid;
  wire                debounce_1_keyStatus_49_payload;
  wire                debounce_1_keyStatus_50_valid;
  wire                debounce_1_keyStatus_50_payload;
  wire                debounce_1_keyStatus_51_valid;
  wire                debounce_1_keyStatus_51_payload;
  wire                debounce_1_keyStatus_52_valid;
  wire                debounce_1_keyStatus_52_payload;
  wire                debounce_1_keyStatus_53_valid;
  wire                debounce_1_keyStatus_53_payload;
  wire                debounce_1_keyStatus_54_valid;
  wire                debounce_1_keyStatus_54_payload;
  wire                debounce_1_keyStatus_55_valid;
  wire                debounce_1_keyStatus_55_payload;
  wire                debounce_1_keyStatus_56_valid;
  wire                debounce_1_keyStatus_56_payload;
  wire                debounce_1_keyStatus_57_valid;
  wire                debounce_1_keyStatus_57_payload;
  wire                debounce_1_keyStatus_58_valid;
  wire                debounce_1_keyStatus_58_payload;
  wire                debounce_1_keyStatus_59_valid;
  wire                debounce_1_keyStatus_59_payload;
  wire                debounce_1_keyStatus_60_valid;
  wire                debounce_1_keyStatus_60_payload;
  wire                debounce_1_keyStatus_61_valid;
  wire                debounce_1_keyStatus_61_payload;
  wire                debounce_1_keyStatus_62_valid;
  wire                debounce_1_keyStatus_62_payload;
  wire                debounce_1_keyStatus_63_valid;
  wire                debounce_1_keyStatus_63_payload;
  wire                debounce_1_keyStatus_64_valid;
  wire                debounce_1_keyStatus_64_payload;
  wire                debounce_1_keyStatus_65_valid;
  wire                debounce_1_keyStatus_65_payload;
  wire                debounce_1_keyStatus_66_valid;
  wire                debounce_1_keyStatus_66_payload;
  wire                debounce_1_keyStatus_67_valid;
  wire                debounce_1_keyStatus_67_payload;
  wire                debounce_1_keyStatus_68_valid;
  wire                debounce_1_keyStatus_68_payload;
  wire                debounce_1_keyStatus_69_valid;
  wire                debounce_1_keyStatus_69_payload;
  wire                debounce_1_keyStatus_70_valid;
  wire                debounce_1_keyStatus_70_payload;
  wire                debounce_1_keyStatus_71_valid;
  wire                debounce_1_keyStatus_71_payload;
  wire                debounce_1_keyStatus_72_valid;
  wire                debounce_1_keyStatus_72_payload;
  wire                debounce_1_keyStatus_73_valid;
  wire                debounce_1_keyStatus_73_payload;
  wire                debounce_1_keyStatus_74_valid;
  wire                debounce_1_keyStatus_74_payload;
  wire                debounce_1_keyStatus_75_valid;
  wire                debounce_1_keyStatus_75_payload;
  wire                debounce_1_keyStatus_76_valid;
  wire                debounce_1_keyStatus_76_payload;
  wire                debounce_1_keyStatus_77_valid;
  wire                debounce_1_keyStatus_77_payload;
  wire                debounce_1_keyStatus_78_valid;
  wire                debounce_1_keyStatus_78_payload;
  wire                debounce_1_keyStatus_79_valid;
  wire                debounce_1_keyStatus_79_payload;
  wire                debounce_1_keyStatus_80_valid;
  wire                debounce_1_keyStatus_80_payload;
  wire                debounce_1_keyStatus_81_valid;
  wire                debounce_1_keyStatus_81_payload;
  wire                debounce_1_keyStatus_82_valid;
  wire                debounce_1_keyStatus_82_payload;
  wire                debounce_1_keyStatus_83_valid;
  wire                debounce_1_keyStatus_83_payload;
  wire                debounce_1_keyStatus_84_valid;
  wire                debounce_1_keyStatus_84_payload;
  wire                debounce_1_keyStatus_85_valid;
  wire                debounce_1_keyStatus_85_payload;
  wire                debounce_1_keyStatus_86_valid;
  wire                debounce_1_keyStatus_86_payload;
  wire                debounce_1_keyStatus_87_valid;
  wire                debounce_1_keyStatus_87_payload;
  wire                debounce_1_keyStatus_88_valid;
  wire                debounce_1_keyStatus_88_payload;
  wire                debounce_1_keyStatus_89_valid;
  wire                debounce_1_keyStatus_89_payload;
  wire                debounce_1_keyStatus_90_valid;
  wire                debounce_1_keyStatus_90_payload;
  wire                debounce_1_keyStatus_91_valid;
  wire                debounce_1_keyStatus_91_payload;
  wire                debounce_1_keyStatus_92_valid;
  wire                debounce_1_keyStatus_92_payload;
  wire                debounce_1_keyStatus_93_valid;
  wire                debounce_1_keyStatus_93_payload;
  wire                debounce_1_keyStatus_94_valid;
  wire                debounce_1_keyStatus_94_payload;
  wire                debounce_1_keyStatus_95_valid;
  wire                debounce_1_keyStatus_95_payload;
  wire                debounce_1_keyStatus_96_valid;
  wire                debounce_1_keyStatus_96_payload;
  wire                debounce_1_keyStatus_97_valid;
  wire                debounce_1_keyStatus_97_payload;
  wire                debounce_1_keyStatus_98_valid;
  wire                debounce_1_keyStatus_98_payload;
  wire                debounce_1_keyStatus_99_valid;
  wire                debounce_1_keyStatus_99_payload;
  wire                debounce_1_keyStatus_100_valid;
  wire                debounce_1_keyStatus_100_payload;
  wire                debounce_1_keyStatus_101_valid;
  wire                debounce_1_keyStatus_101_payload;
  wire                debounce_1_keyStatus_102_valid;
  wire                debounce_1_keyStatus_102_payload;
  wire       [0:0]    _zz_11;
  wire       [12:0]   _zz_12;
  wire       [0:0]    _zz_13;
  wire       [6:0]    _zz_14;
  reg                 clkScan_state;
  reg                 clkScan_stateRise;
  wire                clkScan_counter_willIncrement;
  reg                 clkScan_counter_willClear;
  reg        [12:0]   clkScan_counter_valueNext;
  reg        [12:0]   clkScan_counter_value;
  wire                clkScan_counter_willOverflowIfInc;
  wire                clkScan_counter_willOverflow;
  reg        [7:0]    _zz_2;
  wire                _zz_3;
  reg                 _zz_3_regNext;
  wire                _zz_4;
  reg        [6:0]    _zz_5;
  reg        [6:0]    _zz_6;
  wire                _zz_7;
  wire                _zz_8;

  assign _zz_11 = clkScan_counter_willIncrement;
  assign _zz_12 = {12'd0, _zz_11};
  assign _zz_13 = _zz_4;
  assign _zz_14 = {6'd0, _zz_13};
  scan_key scanK (
    .clock       (clkScan_state          ), //i
    .reset       (_zz_1                  ), //i
    .enabled     (enabled                ), //i
    .COL         (COL[20:0]              ), //i
    .ROW         (scanK_ROW[5:0]         ), //o
    .key_down    (scanK_key_down[102:0]  )  //o
  );
  Debounce debounce_1 (
    .key_down                 (scanK_key_down[102:0]             ), //i
    .keyStatus_0_valid        (debounce_1_keyStatus_0_valid      ), //o
    .keyStatus_0_payload      (debounce_1_keyStatus_0_payload    ), //o
    .keyStatus_1_valid        (debounce_1_keyStatus_1_valid      ), //o
    .keyStatus_1_payload      (debounce_1_keyStatus_1_payload    ), //o
    .keyStatus_2_valid        (debounce_1_keyStatus_2_valid      ), //o
    .keyStatus_2_payload      (debounce_1_keyStatus_2_payload    ), //o
    .keyStatus_3_valid        (debounce_1_keyStatus_3_valid      ), //o
    .keyStatus_3_payload      (debounce_1_keyStatus_3_payload    ), //o
    .keyStatus_4_valid        (debounce_1_keyStatus_4_valid      ), //o
    .keyStatus_4_payload      (debounce_1_keyStatus_4_payload    ), //o
    .keyStatus_5_valid        (debounce_1_keyStatus_5_valid      ), //o
    .keyStatus_5_payload      (debounce_1_keyStatus_5_payload    ), //o
    .keyStatus_6_valid        (debounce_1_keyStatus_6_valid      ), //o
    .keyStatus_6_payload      (debounce_1_keyStatus_6_payload    ), //o
    .keyStatus_7_valid        (debounce_1_keyStatus_7_valid      ), //o
    .keyStatus_7_payload      (debounce_1_keyStatus_7_payload    ), //o
    .keyStatus_8_valid        (debounce_1_keyStatus_8_valid      ), //o
    .keyStatus_8_payload      (debounce_1_keyStatus_8_payload    ), //o
    .keyStatus_9_valid        (debounce_1_keyStatus_9_valid      ), //o
    .keyStatus_9_payload      (debounce_1_keyStatus_9_payload    ), //o
    .keyStatus_10_valid       (debounce_1_keyStatus_10_valid     ), //o
    .keyStatus_10_payload     (debounce_1_keyStatus_10_payload   ), //o
    .keyStatus_11_valid       (debounce_1_keyStatus_11_valid     ), //o
    .keyStatus_11_payload     (debounce_1_keyStatus_11_payload   ), //o
    .keyStatus_12_valid       (debounce_1_keyStatus_12_valid     ), //o
    .keyStatus_12_payload     (debounce_1_keyStatus_12_payload   ), //o
    .keyStatus_13_valid       (debounce_1_keyStatus_13_valid     ), //o
    .keyStatus_13_payload     (debounce_1_keyStatus_13_payload   ), //o
    .keyStatus_14_valid       (debounce_1_keyStatus_14_valid     ), //o
    .keyStatus_14_payload     (debounce_1_keyStatus_14_payload   ), //o
    .keyStatus_15_valid       (debounce_1_keyStatus_15_valid     ), //o
    .keyStatus_15_payload     (debounce_1_keyStatus_15_payload   ), //o
    .keyStatus_16_valid       (debounce_1_keyStatus_16_valid     ), //o
    .keyStatus_16_payload     (debounce_1_keyStatus_16_payload   ), //o
    .keyStatus_17_valid       (debounce_1_keyStatus_17_valid     ), //o
    .keyStatus_17_payload     (debounce_1_keyStatus_17_payload   ), //o
    .keyStatus_18_valid       (debounce_1_keyStatus_18_valid     ), //o
    .keyStatus_18_payload     (debounce_1_keyStatus_18_payload   ), //o
    .keyStatus_19_valid       (debounce_1_keyStatus_19_valid     ), //o
    .keyStatus_19_payload     (debounce_1_keyStatus_19_payload   ), //o
    .keyStatus_20_valid       (debounce_1_keyStatus_20_valid     ), //o
    .keyStatus_20_payload     (debounce_1_keyStatus_20_payload   ), //o
    .keyStatus_21_valid       (debounce_1_keyStatus_21_valid     ), //o
    .keyStatus_21_payload     (debounce_1_keyStatus_21_payload   ), //o
    .keyStatus_22_valid       (debounce_1_keyStatus_22_valid     ), //o
    .keyStatus_22_payload     (debounce_1_keyStatus_22_payload   ), //o
    .keyStatus_23_valid       (debounce_1_keyStatus_23_valid     ), //o
    .keyStatus_23_payload     (debounce_1_keyStatus_23_payload   ), //o
    .keyStatus_24_valid       (debounce_1_keyStatus_24_valid     ), //o
    .keyStatus_24_payload     (debounce_1_keyStatus_24_payload   ), //o
    .keyStatus_25_valid       (debounce_1_keyStatus_25_valid     ), //o
    .keyStatus_25_payload     (debounce_1_keyStatus_25_payload   ), //o
    .keyStatus_26_valid       (debounce_1_keyStatus_26_valid     ), //o
    .keyStatus_26_payload     (debounce_1_keyStatus_26_payload   ), //o
    .keyStatus_27_valid       (debounce_1_keyStatus_27_valid     ), //o
    .keyStatus_27_payload     (debounce_1_keyStatus_27_payload   ), //o
    .keyStatus_28_valid       (debounce_1_keyStatus_28_valid     ), //o
    .keyStatus_28_payload     (debounce_1_keyStatus_28_payload   ), //o
    .keyStatus_29_valid       (debounce_1_keyStatus_29_valid     ), //o
    .keyStatus_29_payload     (debounce_1_keyStatus_29_payload   ), //o
    .keyStatus_30_valid       (debounce_1_keyStatus_30_valid     ), //o
    .keyStatus_30_payload     (debounce_1_keyStatus_30_payload   ), //o
    .keyStatus_31_valid       (debounce_1_keyStatus_31_valid     ), //o
    .keyStatus_31_payload     (debounce_1_keyStatus_31_payload   ), //o
    .keyStatus_32_valid       (debounce_1_keyStatus_32_valid     ), //o
    .keyStatus_32_payload     (debounce_1_keyStatus_32_payload   ), //o
    .keyStatus_33_valid       (debounce_1_keyStatus_33_valid     ), //o
    .keyStatus_33_payload     (debounce_1_keyStatus_33_payload   ), //o
    .keyStatus_34_valid       (debounce_1_keyStatus_34_valid     ), //o
    .keyStatus_34_payload     (debounce_1_keyStatus_34_payload   ), //o
    .keyStatus_35_valid       (debounce_1_keyStatus_35_valid     ), //o
    .keyStatus_35_payload     (debounce_1_keyStatus_35_payload   ), //o
    .keyStatus_36_valid       (debounce_1_keyStatus_36_valid     ), //o
    .keyStatus_36_payload     (debounce_1_keyStatus_36_payload   ), //o
    .keyStatus_37_valid       (debounce_1_keyStatus_37_valid     ), //o
    .keyStatus_37_payload     (debounce_1_keyStatus_37_payload   ), //o
    .keyStatus_38_valid       (debounce_1_keyStatus_38_valid     ), //o
    .keyStatus_38_payload     (debounce_1_keyStatus_38_payload   ), //o
    .keyStatus_39_valid       (debounce_1_keyStatus_39_valid     ), //o
    .keyStatus_39_payload     (debounce_1_keyStatus_39_payload   ), //o
    .keyStatus_40_valid       (debounce_1_keyStatus_40_valid     ), //o
    .keyStatus_40_payload     (debounce_1_keyStatus_40_payload   ), //o
    .keyStatus_41_valid       (debounce_1_keyStatus_41_valid     ), //o
    .keyStatus_41_payload     (debounce_1_keyStatus_41_payload   ), //o
    .keyStatus_42_valid       (debounce_1_keyStatus_42_valid     ), //o
    .keyStatus_42_payload     (debounce_1_keyStatus_42_payload   ), //o
    .keyStatus_43_valid       (debounce_1_keyStatus_43_valid     ), //o
    .keyStatus_43_payload     (debounce_1_keyStatus_43_payload   ), //o
    .keyStatus_44_valid       (debounce_1_keyStatus_44_valid     ), //o
    .keyStatus_44_payload     (debounce_1_keyStatus_44_payload   ), //o
    .keyStatus_45_valid       (debounce_1_keyStatus_45_valid     ), //o
    .keyStatus_45_payload     (debounce_1_keyStatus_45_payload   ), //o
    .keyStatus_46_valid       (debounce_1_keyStatus_46_valid     ), //o
    .keyStatus_46_payload     (debounce_1_keyStatus_46_payload   ), //o
    .keyStatus_47_valid       (debounce_1_keyStatus_47_valid     ), //o
    .keyStatus_47_payload     (debounce_1_keyStatus_47_payload   ), //o
    .keyStatus_48_valid       (debounce_1_keyStatus_48_valid     ), //o
    .keyStatus_48_payload     (debounce_1_keyStatus_48_payload   ), //o
    .keyStatus_49_valid       (debounce_1_keyStatus_49_valid     ), //o
    .keyStatus_49_payload     (debounce_1_keyStatus_49_payload   ), //o
    .keyStatus_50_valid       (debounce_1_keyStatus_50_valid     ), //o
    .keyStatus_50_payload     (debounce_1_keyStatus_50_payload   ), //o
    .keyStatus_51_valid       (debounce_1_keyStatus_51_valid     ), //o
    .keyStatus_51_payload     (debounce_1_keyStatus_51_payload   ), //o
    .keyStatus_52_valid       (debounce_1_keyStatus_52_valid     ), //o
    .keyStatus_52_payload     (debounce_1_keyStatus_52_payload   ), //o
    .keyStatus_53_valid       (debounce_1_keyStatus_53_valid     ), //o
    .keyStatus_53_payload     (debounce_1_keyStatus_53_payload   ), //o
    .keyStatus_54_valid       (debounce_1_keyStatus_54_valid     ), //o
    .keyStatus_54_payload     (debounce_1_keyStatus_54_payload   ), //o
    .keyStatus_55_valid       (debounce_1_keyStatus_55_valid     ), //o
    .keyStatus_55_payload     (debounce_1_keyStatus_55_payload   ), //o
    .keyStatus_56_valid       (debounce_1_keyStatus_56_valid     ), //o
    .keyStatus_56_payload     (debounce_1_keyStatus_56_payload   ), //o
    .keyStatus_57_valid       (debounce_1_keyStatus_57_valid     ), //o
    .keyStatus_57_payload     (debounce_1_keyStatus_57_payload   ), //o
    .keyStatus_58_valid       (debounce_1_keyStatus_58_valid     ), //o
    .keyStatus_58_payload     (debounce_1_keyStatus_58_payload   ), //o
    .keyStatus_59_valid       (debounce_1_keyStatus_59_valid     ), //o
    .keyStatus_59_payload     (debounce_1_keyStatus_59_payload   ), //o
    .keyStatus_60_valid       (debounce_1_keyStatus_60_valid     ), //o
    .keyStatus_60_payload     (debounce_1_keyStatus_60_payload   ), //o
    .keyStatus_61_valid       (debounce_1_keyStatus_61_valid     ), //o
    .keyStatus_61_payload     (debounce_1_keyStatus_61_payload   ), //o
    .keyStatus_62_valid       (debounce_1_keyStatus_62_valid     ), //o
    .keyStatus_62_payload     (debounce_1_keyStatus_62_payload   ), //o
    .keyStatus_63_valid       (debounce_1_keyStatus_63_valid     ), //o
    .keyStatus_63_payload     (debounce_1_keyStatus_63_payload   ), //o
    .keyStatus_64_valid       (debounce_1_keyStatus_64_valid     ), //o
    .keyStatus_64_payload     (debounce_1_keyStatus_64_payload   ), //o
    .keyStatus_65_valid       (debounce_1_keyStatus_65_valid     ), //o
    .keyStatus_65_payload     (debounce_1_keyStatus_65_payload   ), //o
    .keyStatus_66_valid       (debounce_1_keyStatus_66_valid     ), //o
    .keyStatus_66_payload     (debounce_1_keyStatus_66_payload   ), //o
    .keyStatus_67_valid       (debounce_1_keyStatus_67_valid     ), //o
    .keyStatus_67_payload     (debounce_1_keyStatus_67_payload   ), //o
    .keyStatus_68_valid       (debounce_1_keyStatus_68_valid     ), //o
    .keyStatus_68_payload     (debounce_1_keyStatus_68_payload   ), //o
    .keyStatus_69_valid       (debounce_1_keyStatus_69_valid     ), //o
    .keyStatus_69_payload     (debounce_1_keyStatus_69_payload   ), //o
    .keyStatus_70_valid       (debounce_1_keyStatus_70_valid     ), //o
    .keyStatus_70_payload     (debounce_1_keyStatus_70_payload   ), //o
    .keyStatus_71_valid       (debounce_1_keyStatus_71_valid     ), //o
    .keyStatus_71_payload     (debounce_1_keyStatus_71_payload   ), //o
    .keyStatus_72_valid       (debounce_1_keyStatus_72_valid     ), //o
    .keyStatus_72_payload     (debounce_1_keyStatus_72_payload   ), //o
    .keyStatus_73_valid       (debounce_1_keyStatus_73_valid     ), //o
    .keyStatus_73_payload     (debounce_1_keyStatus_73_payload   ), //o
    .keyStatus_74_valid       (debounce_1_keyStatus_74_valid     ), //o
    .keyStatus_74_payload     (debounce_1_keyStatus_74_payload   ), //o
    .keyStatus_75_valid       (debounce_1_keyStatus_75_valid     ), //o
    .keyStatus_75_payload     (debounce_1_keyStatus_75_payload   ), //o
    .keyStatus_76_valid       (debounce_1_keyStatus_76_valid     ), //o
    .keyStatus_76_payload     (debounce_1_keyStatus_76_payload   ), //o
    .keyStatus_77_valid       (debounce_1_keyStatus_77_valid     ), //o
    .keyStatus_77_payload     (debounce_1_keyStatus_77_payload   ), //o
    .keyStatus_78_valid       (debounce_1_keyStatus_78_valid     ), //o
    .keyStatus_78_payload     (debounce_1_keyStatus_78_payload   ), //o
    .keyStatus_79_valid       (debounce_1_keyStatus_79_valid     ), //o
    .keyStatus_79_payload     (debounce_1_keyStatus_79_payload   ), //o
    .keyStatus_80_valid       (debounce_1_keyStatus_80_valid     ), //o
    .keyStatus_80_payload     (debounce_1_keyStatus_80_payload   ), //o
    .keyStatus_81_valid       (debounce_1_keyStatus_81_valid     ), //o
    .keyStatus_81_payload     (debounce_1_keyStatus_81_payload   ), //o
    .keyStatus_82_valid       (debounce_1_keyStatus_82_valid     ), //o
    .keyStatus_82_payload     (debounce_1_keyStatus_82_payload   ), //o
    .keyStatus_83_valid       (debounce_1_keyStatus_83_valid     ), //o
    .keyStatus_83_payload     (debounce_1_keyStatus_83_payload   ), //o
    .keyStatus_84_valid       (debounce_1_keyStatus_84_valid     ), //o
    .keyStatus_84_payload     (debounce_1_keyStatus_84_payload   ), //o
    .keyStatus_85_valid       (debounce_1_keyStatus_85_valid     ), //o
    .keyStatus_85_payload     (debounce_1_keyStatus_85_payload   ), //o
    .keyStatus_86_valid       (debounce_1_keyStatus_86_valid     ), //o
    .keyStatus_86_payload     (debounce_1_keyStatus_86_payload   ), //o
    .keyStatus_87_valid       (debounce_1_keyStatus_87_valid     ), //o
    .keyStatus_87_payload     (debounce_1_keyStatus_87_payload   ), //o
    .keyStatus_88_valid       (debounce_1_keyStatus_88_valid     ), //o
    .keyStatus_88_payload     (debounce_1_keyStatus_88_payload   ), //o
    .keyStatus_89_valid       (debounce_1_keyStatus_89_valid     ), //o
    .keyStatus_89_payload     (debounce_1_keyStatus_89_payload   ), //o
    .keyStatus_90_valid       (debounce_1_keyStatus_90_valid     ), //o
    .keyStatus_90_payload     (debounce_1_keyStatus_90_payload   ), //o
    .keyStatus_91_valid       (debounce_1_keyStatus_91_valid     ), //o
    .keyStatus_91_payload     (debounce_1_keyStatus_91_payload   ), //o
    .keyStatus_92_valid       (debounce_1_keyStatus_92_valid     ), //o
    .keyStatus_92_payload     (debounce_1_keyStatus_92_payload   ), //o
    .keyStatus_93_valid       (debounce_1_keyStatus_93_valid     ), //o
    .keyStatus_93_payload     (debounce_1_keyStatus_93_payload   ), //o
    .keyStatus_94_valid       (debounce_1_keyStatus_94_valid     ), //o
    .keyStatus_94_payload     (debounce_1_keyStatus_94_payload   ), //o
    .keyStatus_95_valid       (debounce_1_keyStatus_95_valid     ), //o
    .keyStatus_95_payload     (debounce_1_keyStatus_95_payload   ), //o
    .keyStatus_96_valid       (debounce_1_keyStatus_96_valid     ), //o
    .keyStatus_96_payload     (debounce_1_keyStatus_96_payload   ), //o
    .keyStatus_97_valid       (debounce_1_keyStatus_97_valid     ), //o
    .keyStatus_97_payload     (debounce_1_keyStatus_97_payload   ), //o
    .keyStatus_98_valid       (debounce_1_keyStatus_98_valid     ), //o
    .keyStatus_98_payload     (debounce_1_keyStatus_98_payload   ), //o
    .keyStatus_99_valid       (debounce_1_keyStatus_99_valid     ), //o
    .keyStatus_99_payload     (debounce_1_keyStatus_99_payload   ), //o
    .keyStatus_100_valid      (debounce_1_keyStatus_100_valid    ), //o
    .keyStatus_100_payload    (debounce_1_keyStatus_100_payload  ), //o
    .keyStatus_101_valid      (debounce_1_keyStatus_101_valid    ), //o
    .keyStatus_101_payload    (debounce_1_keyStatus_101_payload  ), //o
    .keyStatus_102_valid      (debounce_1_keyStatus_102_valid    ), //o
    .keyStatus_102_payload    (debounce_1_keyStatus_102_payload  ), //o
    .CLK_50                   (CLK_50                            ), //i
    ._zz_3                    (_zz_1                             )  //i
  );
  always @(*) begin
    case(_zz_6)
      7'b0000000 : begin
        _zz_9 = keyStatus_0_valid;
        _zz_10 = keyStatus_0_payload;
      end
      7'b0000001 : begin
        _zz_9 = keyStatus_1_valid;
        _zz_10 = keyStatus_1_payload;
      end
      7'b0000010 : begin
        _zz_9 = keyStatus_2_valid;
        _zz_10 = keyStatus_2_payload;
      end
      7'b0000011 : begin
        _zz_9 = keyStatus_3_valid;
        _zz_10 = keyStatus_3_payload;
      end
      7'b0000100 : begin
        _zz_9 = keyStatus_4_valid;
        _zz_10 = keyStatus_4_payload;
      end
      7'b0000101 : begin
        _zz_9 = keyStatus_5_valid;
        _zz_10 = keyStatus_5_payload;
      end
      7'b0000110 : begin
        _zz_9 = keyStatus_6_valid;
        _zz_10 = keyStatus_6_payload;
      end
      7'b0000111 : begin
        _zz_9 = keyStatus_7_valid;
        _zz_10 = keyStatus_7_payload;
      end
      7'b0001000 : begin
        _zz_9 = keyStatus_8_valid;
        _zz_10 = keyStatus_8_payload;
      end
      7'b0001001 : begin
        _zz_9 = keyStatus_9_valid;
        _zz_10 = keyStatus_9_payload;
      end
      7'b0001010 : begin
        _zz_9 = keyStatus_10_valid;
        _zz_10 = keyStatus_10_payload;
      end
      7'b0001011 : begin
        _zz_9 = keyStatus_11_valid;
        _zz_10 = keyStatus_11_payload;
      end
      7'b0001100 : begin
        _zz_9 = keyStatus_12_valid;
        _zz_10 = keyStatus_12_payload;
      end
      7'b0001101 : begin
        _zz_9 = keyStatus_13_valid;
        _zz_10 = keyStatus_13_payload;
      end
      7'b0001110 : begin
        _zz_9 = keyStatus_14_valid;
        _zz_10 = keyStatus_14_payload;
      end
      7'b0001111 : begin
        _zz_9 = keyStatus_15_valid;
        _zz_10 = keyStatus_15_payload;
      end
      7'b0010000 : begin
        _zz_9 = keyStatus_16_valid;
        _zz_10 = keyStatus_16_payload;
      end
      7'b0010001 : begin
        _zz_9 = keyStatus_17_valid;
        _zz_10 = keyStatus_17_payload;
      end
      7'b0010010 : begin
        _zz_9 = keyStatus_18_valid;
        _zz_10 = keyStatus_18_payload;
      end
      7'b0010011 : begin
        _zz_9 = keyStatus_19_valid;
        _zz_10 = keyStatus_19_payload;
      end
      7'b0010100 : begin
        _zz_9 = keyStatus_20_valid;
        _zz_10 = keyStatus_20_payload;
      end
      7'b0010101 : begin
        _zz_9 = keyStatus_21_valid;
        _zz_10 = keyStatus_21_payload;
      end
      7'b0010110 : begin
        _zz_9 = keyStatus_22_valid;
        _zz_10 = keyStatus_22_payload;
      end
      7'b0010111 : begin
        _zz_9 = keyStatus_23_valid;
        _zz_10 = keyStatus_23_payload;
      end
      7'b0011000 : begin
        _zz_9 = keyStatus_24_valid;
        _zz_10 = keyStatus_24_payload;
      end
      7'b0011001 : begin
        _zz_9 = keyStatus_25_valid;
        _zz_10 = keyStatus_25_payload;
      end
      7'b0011010 : begin
        _zz_9 = keyStatus_26_valid;
        _zz_10 = keyStatus_26_payload;
      end
      7'b0011011 : begin
        _zz_9 = keyStatus_27_valid;
        _zz_10 = keyStatus_27_payload;
      end
      7'b0011100 : begin
        _zz_9 = keyStatus_28_valid;
        _zz_10 = keyStatus_28_payload;
      end
      7'b0011101 : begin
        _zz_9 = keyStatus_29_valid;
        _zz_10 = keyStatus_29_payload;
      end
      7'b0011110 : begin
        _zz_9 = keyStatus_30_valid;
        _zz_10 = keyStatus_30_payload;
      end
      7'b0011111 : begin
        _zz_9 = keyStatus_31_valid;
        _zz_10 = keyStatus_31_payload;
      end
      7'b0100000 : begin
        _zz_9 = keyStatus_32_valid;
        _zz_10 = keyStatus_32_payload;
      end
      7'b0100001 : begin
        _zz_9 = keyStatus_33_valid;
        _zz_10 = keyStatus_33_payload;
      end
      7'b0100010 : begin
        _zz_9 = keyStatus_34_valid;
        _zz_10 = keyStatus_34_payload;
      end
      7'b0100011 : begin
        _zz_9 = keyStatus_35_valid;
        _zz_10 = keyStatus_35_payload;
      end
      7'b0100100 : begin
        _zz_9 = keyStatus_36_valid;
        _zz_10 = keyStatus_36_payload;
      end
      7'b0100101 : begin
        _zz_9 = keyStatus_37_valid;
        _zz_10 = keyStatus_37_payload;
      end
      7'b0100110 : begin
        _zz_9 = keyStatus_38_valid;
        _zz_10 = keyStatus_38_payload;
      end
      7'b0100111 : begin
        _zz_9 = keyStatus_39_valid;
        _zz_10 = keyStatus_39_payload;
      end
      7'b0101000 : begin
        _zz_9 = keyStatus_40_valid;
        _zz_10 = keyStatus_40_payload;
      end
      7'b0101001 : begin
        _zz_9 = keyStatus_41_valid;
        _zz_10 = keyStatus_41_payload;
      end
      7'b0101010 : begin
        _zz_9 = keyStatus_42_valid;
        _zz_10 = keyStatus_42_payload;
      end
      7'b0101011 : begin
        _zz_9 = keyStatus_43_valid;
        _zz_10 = keyStatus_43_payload;
      end
      7'b0101100 : begin
        _zz_9 = keyStatus_44_valid;
        _zz_10 = keyStatus_44_payload;
      end
      7'b0101101 : begin
        _zz_9 = keyStatus_45_valid;
        _zz_10 = keyStatus_45_payload;
      end
      7'b0101110 : begin
        _zz_9 = keyStatus_46_valid;
        _zz_10 = keyStatus_46_payload;
      end
      7'b0101111 : begin
        _zz_9 = keyStatus_47_valid;
        _zz_10 = keyStatus_47_payload;
      end
      7'b0110000 : begin
        _zz_9 = keyStatus_48_valid;
        _zz_10 = keyStatus_48_payload;
      end
      7'b0110001 : begin
        _zz_9 = keyStatus_49_valid;
        _zz_10 = keyStatus_49_payload;
      end
      7'b0110010 : begin
        _zz_9 = keyStatus_50_valid;
        _zz_10 = keyStatus_50_payload;
      end
      7'b0110011 : begin
        _zz_9 = keyStatus_51_valid;
        _zz_10 = keyStatus_51_payload;
      end
      7'b0110100 : begin
        _zz_9 = keyStatus_52_valid;
        _zz_10 = keyStatus_52_payload;
      end
      7'b0110101 : begin
        _zz_9 = keyStatus_53_valid;
        _zz_10 = keyStatus_53_payload;
      end
      7'b0110110 : begin
        _zz_9 = keyStatus_54_valid;
        _zz_10 = keyStatus_54_payload;
      end
      7'b0110111 : begin
        _zz_9 = keyStatus_55_valid;
        _zz_10 = keyStatus_55_payload;
      end
      7'b0111000 : begin
        _zz_9 = keyStatus_56_valid;
        _zz_10 = keyStatus_56_payload;
      end
      7'b0111001 : begin
        _zz_9 = keyStatus_57_valid;
        _zz_10 = keyStatus_57_payload;
      end
      7'b0111010 : begin
        _zz_9 = keyStatus_58_valid;
        _zz_10 = keyStatus_58_payload;
      end
      7'b0111011 : begin
        _zz_9 = keyStatus_59_valid;
        _zz_10 = keyStatus_59_payload;
      end
      7'b0111100 : begin
        _zz_9 = keyStatus_60_valid;
        _zz_10 = keyStatus_60_payload;
      end
      7'b0111101 : begin
        _zz_9 = keyStatus_61_valid;
        _zz_10 = keyStatus_61_payload;
      end
      7'b0111110 : begin
        _zz_9 = keyStatus_62_valid;
        _zz_10 = keyStatus_62_payload;
      end
      7'b0111111 : begin
        _zz_9 = keyStatus_63_valid;
        _zz_10 = keyStatus_63_payload;
      end
      7'b1000000 : begin
        _zz_9 = keyStatus_64_valid;
        _zz_10 = keyStatus_64_payload;
      end
      7'b1000001 : begin
        _zz_9 = keyStatus_65_valid;
        _zz_10 = keyStatus_65_payload;
      end
      7'b1000010 : begin
        _zz_9 = keyStatus_66_valid;
        _zz_10 = keyStatus_66_payload;
      end
      7'b1000011 : begin
        _zz_9 = keyStatus_67_valid;
        _zz_10 = keyStatus_67_payload;
      end
      7'b1000100 : begin
        _zz_9 = keyStatus_68_valid;
        _zz_10 = keyStatus_68_payload;
      end
      7'b1000101 : begin
        _zz_9 = keyStatus_69_valid;
        _zz_10 = keyStatus_69_payload;
      end
      7'b1000110 : begin
        _zz_9 = keyStatus_70_valid;
        _zz_10 = keyStatus_70_payload;
      end
      7'b1000111 : begin
        _zz_9 = keyStatus_71_valid;
        _zz_10 = keyStatus_71_payload;
      end
      7'b1001000 : begin
        _zz_9 = keyStatus_72_valid;
        _zz_10 = keyStatus_72_payload;
      end
      7'b1001001 : begin
        _zz_9 = keyStatus_73_valid;
        _zz_10 = keyStatus_73_payload;
      end
      7'b1001010 : begin
        _zz_9 = keyStatus_74_valid;
        _zz_10 = keyStatus_74_payload;
      end
      7'b1001011 : begin
        _zz_9 = keyStatus_75_valid;
        _zz_10 = keyStatus_75_payload;
      end
      7'b1001100 : begin
        _zz_9 = keyStatus_76_valid;
        _zz_10 = keyStatus_76_payload;
      end
      7'b1001101 : begin
        _zz_9 = keyStatus_77_valid;
        _zz_10 = keyStatus_77_payload;
      end
      7'b1001110 : begin
        _zz_9 = keyStatus_78_valid;
        _zz_10 = keyStatus_78_payload;
      end
      7'b1001111 : begin
        _zz_9 = keyStatus_79_valid;
        _zz_10 = keyStatus_79_payload;
      end
      7'b1010000 : begin
        _zz_9 = keyStatus_80_valid;
        _zz_10 = keyStatus_80_payload;
      end
      7'b1010001 : begin
        _zz_9 = keyStatus_81_valid;
        _zz_10 = keyStatus_81_payload;
      end
      7'b1010010 : begin
        _zz_9 = keyStatus_82_valid;
        _zz_10 = keyStatus_82_payload;
      end
      7'b1010011 : begin
        _zz_9 = keyStatus_83_valid;
        _zz_10 = keyStatus_83_payload;
      end
      7'b1010100 : begin
        _zz_9 = keyStatus_84_valid;
        _zz_10 = keyStatus_84_payload;
      end
      7'b1010101 : begin
        _zz_9 = keyStatus_85_valid;
        _zz_10 = keyStatus_85_payload;
      end
      7'b1010110 : begin
        _zz_9 = keyStatus_86_valid;
        _zz_10 = keyStatus_86_payload;
      end
      7'b1010111 : begin
        _zz_9 = keyStatus_87_valid;
        _zz_10 = keyStatus_87_payload;
      end
      7'b1011000 : begin
        _zz_9 = keyStatus_88_valid;
        _zz_10 = keyStatus_88_payload;
      end
      7'b1011001 : begin
        _zz_9 = keyStatus_89_valid;
        _zz_10 = keyStatus_89_payload;
      end
      7'b1011010 : begin
        _zz_9 = keyStatus_90_valid;
        _zz_10 = keyStatus_90_payload;
      end
      7'b1011011 : begin
        _zz_9 = keyStatus_91_valid;
        _zz_10 = keyStatus_91_payload;
      end
      7'b1011100 : begin
        _zz_9 = keyStatus_92_valid;
        _zz_10 = keyStatus_92_payload;
      end
      7'b1011101 : begin
        _zz_9 = keyStatus_93_valid;
        _zz_10 = keyStatus_93_payload;
      end
      7'b1011110 : begin
        _zz_9 = keyStatus_94_valid;
        _zz_10 = keyStatus_94_payload;
      end
      7'b1011111 : begin
        _zz_9 = keyStatus_95_valid;
        _zz_10 = keyStatus_95_payload;
      end
      7'b1100000 : begin
        _zz_9 = keyStatus_96_valid;
        _zz_10 = keyStatus_96_payload;
      end
      7'b1100001 : begin
        _zz_9 = keyStatus_97_valid;
        _zz_10 = keyStatus_97_payload;
      end
      7'b1100010 : begin
        _zz_9 = keyStatus_98_valid;
        _zz_10 = keyStatus_98_payload;
      end
      7'b1100011 : begin
        _zz_9 = keyStatus_99_valid;
        _zz_10 = keyStatus_99_payload;
      end
      7'b1100100 : begin
        _zz_9 = keyStatus_100_valid;
        _zz_10 = keyStatus_100_payload;
      end
      7'b1100101 : begin
        _zz_9 = keyStatus_101_valid;
        _zz_10 = keyStatus_101_payload;
      end
      default : begin
        _zz_9 = keyStatus_102_valid;
        _zz_10 = keyStatus_102_payload;
      end
    endcase
  end

  always @ (*) begin
    clkScan_stateRise = 1'b0;
    if(clkScan_counter_willOverflow)begin
      clkScan_stateRise = (! clkScan_state);
    end
    if(clkScan_state)begin
      clkScan_stateRise = 1'b0;
    end
  end

  always @ (*) begin
    clkScan_counter_willClear = 1'b0;
    if(clkScan_state)begin
      clkScan_counter_willClear = 1'b1;
    end
  end

  assign clkScan_counter_willOverflowIfInc = (clkScan_counter_value == 13'h1045);
  assign clkScan_counter_willOverflow = (clkScan_counter_willOverflowIfInc && clkScan_counter_willIncrement);
  always @ (*) begin
    if(clkScan_counter_willOverflow)begin
      clkScan_counter_valueNext = 13'h0;
    end else begin
      clkScan_counter_valueNext = (clkScan_counter_value + _zz_12);
    end
    if(clkScan_counter_willClear)begin
      clkScan_counter_valueNext = 13'h0;
    end
  end

  assign clkScan_counter_willIncrement = 1'b1;
  assign ROW = scanK_ROW;
  assign keyStatus_0_valid = debounce_1_keyStatus_0_valid;
  assign keyStatus_0_payload = debounce_1_keyStatus_0_payload;
  assign keyStatus_1_valid = debounce_1_keyStatus_1_valid;
  assign keyStatus_1_payload = debounce_1_keyStatus_1_payload;
  assign keyStatus_2_valid = debounce_1_keyStatus_2_valid;
  assign keyStatus_2_payload = debounce_1_keyStatus_2_payload;
  assign keyStatus_3_valid = debounce_1_keyStatus_3_valid;
  assign keyStatus_3_payload = debounce_1_keyStatus_3_payload;
  assign keyStatus_4_valid = debounce_1_keyStatus_4_valid;
  assign keyStatus_4_payload = debounce_1_keyStatus_4_payload;
  assign keyStatus_5_valid = debounce_1_keyStatus_5_valid;
  assign keyStatus_5_payload = debounce_1_keyStatus_5_payload;
  assign keyStatus_6_valid = debounce_1_keyStatus_6_valid;
  assign keyStatus_6_payload = debounce_1_keyStatus_6_payload;
  assign keyStatus_7_valid = debounce_1_keyStatus_7_valid;
  assign keyStatus_7_payload = debounce_1_keyStatus_7_payload;
  assign keyStatus_8_valid = debounce_1_keyStatus_8_valid;
  assign keyStatus_8_payload = debounce_1_keyStatus_8_payload;
  assign keyStatus_9_valid = debounce_1_keyStatus_9_valid;
  assign keyStatus_9_payload = debounce_1_keyStatus_9_payload;
  assign keyStatus_10_valid = debounce_1_keyStatus_10_valid;
  assign keyStatus_10_payload = debounce_1_keyStatus_10_payload;
  assign keyStatus_11_valid = debounce_1_keyStatus_11_valid;
  assign keyStatus_11_payload = debounce_1_keyStatus_11_payload;
  assign keyStatus_12_valid = debounce_1_keyStatus_12_valid;
  assign keyStatus_12_payload = debounce_1_keyStatus_12_payload;
  assign keyStatus_13_valid = debounce_1_keyStatus_13_valid;
  assign keyStatus_13_payload = debounce_1_keyStatus_13_payload;
  assign keyStatus_14_valid = debounce_1_keyStatus_14_valid;
  assign keyStatus_14_payload = debounce_1_keyStatus_14_payload;
  assign keyStatus_15_valid = debounce_1_keyStatus_15_valid;
  assign keyStatus_15_payload = debounce_1_keyStatus_15_payload;
  assign keyStatus_16_valid = debounce_1_keyStatus_16_valid;
  assign keyStatus_16_payload = debounce_1_keyStatus_16_payload;
  assign keyStatus_17_valid = debounce_1_keyStatus_17_valid;
  assign keyStatus_17_payload = debounce_1_keyStatus_17_payload;
  assign keyStatus_18_valid = debounce_1_keyStatus_18_valid;
  assign keyStatus_18_payload = debounce_1_keyStatus_18_payload;
  assign keyStatus_19_valid = debounce_1_keyStatus_19_valid;
  assign keyStatus_19_payload = debounce_1_keyStatus_19_payload;
  assign keyStatus_20_valid = debounce_1_keyStatus_20_valid;
  assign keyStatus_20_payload = debounce_1_keyStatus_20_payload;
  assign keyStatus_21_valid = debounce_1_keyStatus_21_valid;
  assign keyStatus_21_payload = debounce_1_keyStatus_21_payload;
  assign keyStatus_22_valid = debounce_1_keyStatus_22_valid;
  assign keyStatus_22_payload = debounce_1_keyStatus_22_payload;
  assign keyStatus_23_valid = debounce_1_keyStatus_23_valid;
  assign keyStatus_23_payload = debounce_1_keyStatus_23_payload;
  assign keyStatus_24_valid = debounce_1_keyStatus_24_valid;
  assign keyStatus_24_payload = debounce_1_keyStatus_24_payload;
  assign keyStatus_25_valid = debounce_1_keyStatus_25_valid;
  assign keyStatus_25_payload = debounce_1_keyStatus_25_payload;
  assign keyStatus_26_valid = debounce_1_keyStatus_26_valid;
  assign keyStatus_26_payload = debounce_1_keyStatus_26_payload;
  assign keyStatus_27_valid = debounce_1_keyStatus_27_valid;
  assign keyStatus_27_payload = debounce_1_keyStatus_27_payload;
  assign keyStatus_28_valid = debounce_1_keyStatus_28_valid;
  assign keyStatus_28_payload = debounce_1_keyStatus_28_payload;
  assign keyStatus_29_valid = debounce_1_keyStatus_29_valid;
  assign keyStatus_29_payload = debounce_1_keyStatus_29_payload;
  assign keyStatus_30_valid = debounce_1_keyStatus_30_valid;
  assign keyStatus_30_payload = debounce_1_keyStatus_30_payload;
  assign keyStatus_31_valid = debounce_1_keyStatus_31_valid;
  assign keyStatus_31_payload = debounce_1_keyStatus_31_payload;
  assign keyStatus_32_valid = debounce_1_keyStatus_32_valid;
  assign keyStatus_32_payload = debounce_1_keyStatus_32_payload;
  assign keyStatus_33_valid = debounce_1_keyStatus_33_valid;
  assign keyStatus_33_payload = debounce_1_keyStatus_33_payload;
  assign keyStatus_34_valid = debounce_1_keyStatus_34_valid;
  assign keyStatus_34_payload = debounce_1_keyStatus_34_payload;
  assign keyStatus_35_valid = debounce_1_keyStatus_35_valid;
  assign keyStatus_35_payload = debounce_1_keyStatus_35_payload;
  assign keyStatus_36_valid = debounce_1_keyStatus_36_valid;
  assign keyStatus_36_payload = debounce_1_keyStatus_36_payload;
  assign keyStatus_37_valid = debounce_1_keyStatus_37_valid;
  assign keyStatus_37_payload = debounce_1_keyStatus_37_payload;
  assign keyStatus_38_valid = debounce_1_keyStatus_38_valid;
  assign keyStatus_38_payload = debounce_1_keyStatus_38_payload;
  assign keyStatus_39_valid = debounce_1_keyStatus_39_valid;
  assign keyStatus_39_payload = debounce_1_keyStatus_39_payload;
  assign keyStatus_40_valid = debounce_1_keyStatus_40_valid;
  assign keyStatus_40_payload = debounce_1_keyStatus_40_payload;
  assign keyStatus_41_valid = debounce_1_keyStatus_41_valid;
  assign keyStatus_41_payload = debounce_1_keyStatus_41_payload;
  assign keyStatus_42_valid = debounce_1_keyStatus_42_valid;
  assign keyStatus_42_payload = debounce_1_keyStatus_42_payload;
  assign keyStatus_43_valid = debounce_1_keyStatus_43_valid;
  assign keyStatus_43_payload = debounce_1_keyStatus_43_payload;
  assign keyStatus_44_valid = debounce_1_keyStatus_44_valid;
  assign keyStatus_44_payload = debounce_1_keyStatus_44_payload;
  assign keyStatus_45_valid = debounce_1_keyStatus_45_valid;
  assign keyStatus_45_payload = debounce_1_keyStatus_45_payload;
  assign keyStatus_46_valid = debounce_1_keyStatus_46_valid;
  assign keyStatus_46_payload = debounce_1_keyStatus_46_payload;
  assign keyStatus_47_valid = debounce_1_keyStatus_47_valid;
  assign keyStatus_47_payload = debounce_1_keyStatus_47_payload;
  assign keyStatus_48_valid = debounce_1_keyStatus_48_valid;
  assign keyStatus_48_payload = debounce_1_keyStatus_48_payload;
  assign keyStatus_49_valid = debounce_1_keyStatus_49_valid;
  assign keyStatus_49_payload = debounce_1_keyStatus_49_payload;
  assign keyStatus_50_valid = debounce_1_keyStatus_50_valid;
  assign keyStatus_50_payload = debounce_1_keyStatus_50_payload;
  assign keyStatus_51_valid = debounce_1_keyStatus_51_valid;
  assign keyStatus_51_payload = debounce_1_keyStatus_51_payload;
  assign keyStatus_52_valid = debounce_1_keyStatus_52_valid;
  assign keyStatus_52_payload = debounce_1_keyStatus_52_payload;
  assign keyStatus_53_valid = debounce_1_keyStatus_53_valid;
  assign keyStatus_53_payload = debounce_1_keyStatus_53_payload;
  assign keyStatus_54_valid = debounce_1_keyStatus_54_valid;
  assign keyStatus_54_payload = debounce_1_keyStatus_54_payload;
  assign keyStatus_55_valid = debounce_1_keyStatus_55_valid;
  assign keyStatus_55_payload = debounce_1_keyStatus_55_payload;
  assign keyStatus_56_valid = debounce_1_keyStatus_56_valid;
  assign keyStatus_56_payload = debounce_1_keyStatus_56_payload;
  assign keyStatus_57_valid = debounce_1_keyStatus_57_valid;
  assign keyStatus_57_payload = debounce_1_keyStatus_57_payload;
  assign keyStatus_58_valid = debounce_1_keyStatus_58_valid;
  assign keyStatus_58_payload = debounce_1_keyStatus_58_payload;
  assign keyStatus_59_valid = debounce_1_keyStatus_59_valid;
  assign keyStatus_59_payload = debounce_1_keyStatus_59_payload;
  assign keyStatus_60_valid = debounce_1_keyStatus_60_valid;
  assign keyStatus_60_payload = debounce_1_keyStatus_60_payload;
  assign keyStatus_61_valid = debounce_1_keyStatus_61_valid;
  assign keyStatus_61_payload = debounce_1_keyStatus_61_payload;
  assign keyStatus_62_valid = debounce_1_keyStatus_62_valid;
  assign keyStatus_62_payload = debounce_1_keyStatus_62_payload;
  assign keyStatus_63_valid = debounce_1_keyStatus_63_valid;
  assign keyStatus_63_payload = debounce_1_keyStatus_63_payload;
  assign keyStatus_64_valid = debounce_1_keyStatus_64_valid;
  assign keyStatus_64_payload = debounce_1_keyStatus_64_payload;
  assign keyStatus_65_valid = debounce_1_keyStatus_65_valid;
  assign keyStatus_65_payload = debounce_1_keyStatus_65_payload;
  assign keyStatus_66_valid = debounce_1_keyStatus_66_valid;
  assign keyStatus_66_payload = debounce_1_keyStatus_66_payload;
  assign keyStatus_67_valid = debounce_1_keyStatus_67_valid;
  assign keyStatus_67_payload = debounce_1_keyStatus_67_payload;
  assign keyStatus_68_valid = debounce_1_keyStatus_68_valid;
  assign keyStatus_68_payload = debounce_1_keyStatus_68_payload;
  assign keyStatus_69_valid = debounce_1_keyStatus_69_valid;
  assign keyStatus_69_payload = debounce_1_keyStatus_69_payload;
  assign keyStatus_70_valid = debounce_1_keyStatus_70_valid;
  assign keyStatus_70_payload = debounce_1_keyStatus_70_payload;
  assign keyStatus_71_valid = debounce_1_keyStatus_71_valid;
  assign keyStatus_71_payload = debounce_1_keyStatus_71_payload;
  assign keyStatus_72_valid = debounce_1_keyStatus_72_valid;
  assign keyStatus_72_payload = debounce_1_keyStatus_72_payload;
  assign keyStatus_73_valid = debounce_1_keyStatus_73_valid;
  assign keyStatus_73_payload = debounce_1_keyStatus_73_payload;
  assign keyStatus_74_valid = debounce_1_keyStatus_74_valid;
  assign keyStatus_74_payload = debounce_1_keyStatus_74_payload;
  assign keyStatus_75_valid = debounce_1_keyStatus_75_valid;
  assign keyStatus_75_payload = debounce_1_keyStatus_75_payload;
  assign keyStatus_76_valid = debounce_1_keyStatus_76_valid;
  assign keyStatus_76_payload = debounce_1_keyStatus_76_payload;
  assign keyStatus_77_valid = debounce_1_keyStatus_77_valid;
  assign keyStatus_77_payload = debounce_1_keyStatus_77_payload;
  assign keyStatus_78_valid = debounce_1_keyStatus_78_valid;
  assign keyStatus_78_payload = debounce_1_keyStatus_78_payload;
  assign keyStatus_79_valid = debounce_1_keyStatus_79_valid;
  assign keyStatus_79_payload = debounce_1_keyStatus_79_payload;
  assign keyStatus_80_valid = debounce_1_keyStatus_80_valid;
  assign keyStatus_80_payload = debounce_1_keyStatus_80_payload;
  assign keyStatus_81_valid = debounce_1_keyStatus_81_valid;
  assign keyStatus_81_payload = debounce_1_keyStatus_81_payload;
  assign keyStatus_82_valid = debounce_1_keyStatus_82_valid;
  assign keyStatus_82_payload = debounce_1_keyStatus_82_payload;
  assign keyStatus_83_valid = debounce_1_keyStatus_83_valid;
  assign keyStatus_83_payload = debounce_1_keyStatus_83_payload;
  assign keyStatus_84_valid = debounce_1_keyStatus_84_valid;
  assign keyStatus_84_payload = debounce_1_keyStatus_84_payload;
  assign keyStatus_85_valid = debounce_1_keyStatus_85_valid;
  assign keyStatus_85_payload = debounce_1_keyStatus_85_payload;
  assign keyStatus_86_valid = debounce_1_keyStatus_86_valid;
  assign keyStatus_86_payload = debounce_1_keyStatus_86_payload;
  assign keyStatus_87_valid = debounce_1_keyStatus_87_valid;
  assign keyStatus_87_payload = debounce_1_keyStatus_87_payload;
  assign keyStatus_88_valid = debounce_1_keyStatus_88_valid;
  assign keyStatus_88_payload = debounce_1_keyStatus_88_payload;
  assign keyStatus_89_valid = debounce_1_keyStatus_89_valid;
  assign keyStatus_89_payload = debounce_1_keyStatus_89_payload;
  assign keyStatus_90_valid = debounce_1_keyStatus_90_valid;
  assign keyStatus_90_payload = debounce_1_keyStatus_90_payload;
  assign keyStatus_91_valid = debounce_1_keyStatus_91_valid;
  assign keyStatus_91_payload = debounce_1_keyStatus_91_payload;
  assign keyStatus_92_valid = debounce_1_keyStatus_92_valid;
  assign keyStatus_92_payload = debounce_1_keyStatus_92_payload;
  assign keyStatus_93_valid = debounce_1_keyStatus_93_valid;
  assign keyStatus_93_payload = debounce_1_keyStatus_93_payload;
  assign keyStatus_94_valid = debounce_1_keyStatus_94_valid;
  assign keyStatus_94_payload = debounce_1_keyStatus_94_payload;
  assign keyStatus_95_valid = debounce_1_keyStatus_95_valid;
  assign keyStatus_95_payload = debounce_1_keyStatus_95_payload;
  assign keyStatus_96_valid = debounce_1_keyStatus_96_valid;
  assign keyStatus_96_payload = debounce_1_keyStatus_96_payload;
  assign keyStatus_97_valid = debounce_1_keyStatus_97_valid;
  assign keyStatus_97_payload = debounce_1_keyStatus_97_payload;
  assign keyStatus_98_valid = debounce_1_keyStatus_98_valid;
  assign keyStatus_98_payload = debounce_1_keyStatus_98_payload;
  assign keyStatus_99_valid = debounce_1_keyStatus_99_valid;
  assign keyStatus_99_payload = debounce_1_keyStatus_99_payload;
  assign keyStatus_100_valid = debounce_1_keyStatus_100_valid;
  assign keyStatus_100_payload = debounce_1_keyStatus_100_payload;
  assign keyStatus_101_valid = debounce_1_keyStatus_101_valid;
  assign keyStatus_101_payload = debounce_1_keyStatus_101_payload;
  assign keyStatus_102_valid = debounce_1_keyStatus_102_valid;
  assign keyStatus_102_payload = debounce_1_keyStatus_102_payload;
  assign _zz_3 = (_zz_2 == 8'hf1);
  assign _zz_7 = (_zz_6 == 7'h66);
  assign _zz_8 = (_zz_7 && _zz_4);
  always @ (*) begin
    if(_zz_8)begin
      _zz_5 = 7'h0;
    end else begin
      _zz_5 = (_zz_6 + _zz_14);
    end
    if(1'b0)begin
      _zz_5 = 7'h0;
    end
  end

  assign _zz_4 = 1'b1;
  assign scanIdx_valid = _zz_9;
  assign scanIdx_payload = {_zz_10,_zz_6};
  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      clkScan_state <= 1'b0;
      clkScan_counter_value <= 13'h0;
      _zz_2 <= 8'h0;
      _zz_3_regNext <= 1'b0;
    end else begin
      clkScan_counter_value <= clkScan_counter_valueNext;
      if(clkScan_counter_willOverflow)begin
        clkScan_state <= 1'b1;
      end
      if(clkScan_state)begin
        clkScan_state <= 1'b0;
      end
      _zz_2 <= (_zz_2 + 8'h01);
      if(_zz_3)begin
        _zz_2 <= 8'h0;
      end
      _zz_3_regNext <= _zz_3;
    end
  end

  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      _zz_6 <= 7'h0;
    end else begin
      if(_zz_3_regNext) begin
        _zz_6 <= _zz_5;
      end
    end
  end


endmodule

module BufferCC_2 (
  input               io_dataIn,
  output              io_dataOut,
  input               CLK_50,
  input               _zz_1
);
  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module ResetController (
  input               io_clock,
  input               io_externalReset,
  output              io_globalReset
);
  wire       [0:0]    _zz_14;
  wire       [15:0]   _zz_15;
  wire       [0:0]    _zz_16;
  wire       [27:0]   _zz_17;
  reg                 _zz_1;
  reg        [15:0]   _zz_2;
  reg        [15:0]   _zz_3 = 16'h0;
  wire                _zz_4;
  wire                _zz_5;
  reg                 _zz_6 = 1'b1;
  reg                 _zz_7;
  reg                 _zz_8;
  reg        [27:0]   _zz_9;
  reg        [27:0]   _zz_10 = 28'h0;
  wire                _zz_11;
  wire                _zz_12;
  reg                 io_externalReset_regNext = 1'b0;
  reg                 _zz_13;

  assign _zz_14 = _zz_1;
  assign _zz_15 = {15'd0, _zz_14};
  assign _zz_16 = _zz_7;
  assign _zz_17 = {27'd0, _zz_16};
  always @ (*) begin
    _zz_1 = 1'b0;
    if(_zz_6)begin
      _zz_1 = 1'b1;
    end
  end

  assign _zz_4 = (_zz_3 == 16'hc34f);
  assign _zz_5 = (_zz_4 && _zz_1);
  always @ (*) begin
    if(_zz_5)begin
      _zz_2 = 16'h0;
    end else begin
      _zz_2 = (_zz_3 + _zz_15);
    end
    if(1'b0)begin
      _zz_2 = 16'h0;
    end
  end

  always @ (*) begin
    _zz_7 = 1'b0;
    if(io_externalReset)begin
      _zz_7 = 1'b1;
    end
  end

  always @ (*) begin
    _zz_8 = 1'b0;
    if((io_externalReset && (! io_externalReset_regNext)))begin
      _zz_8 = 1'b1;
    end
  end

  assign _zz_11 = (_zz_10 == 28'h8f0d17f);
  assign _zz_12 = (_zz_11 && _zz_7);
  always @ (*) begin
    if(_zz_12)begin
      _zz_9 = 28'h0;
    end else begin
      _zz_9 = (_zz_10 + _zz_17);
    end
    if(_zz_8)begin
      _zz_9 = 28'h0;
    end
  end

  assign io_globalReset = _zz_13;
  always @ (posedge io_clock) begin
    _zz_3 <= _zz_2;
    if(_zz_4)begin
      _zz_6 <= 1'b0;
    end
    _zz_10 <= _zz_9;
    io_externalReset_regNext <= io_externalReset;
  end

  always @ (posedge io_clock) begin
    _zz_13 <= (_zz_6 || _zz_12);
  end


endmodule

module UartCtrl (
  input      [2:0]    io_config_frame_dataLength,
  input      `UartStopType_defaultEncoding_type io_config_frame_stop,
  input      `UartParityType_defaultEncoding_type io_config_frame_parity,
  input      [19:0]   io_config_clockDivider,
  input               io_write_valid,
  output reg          io_write_ready,
  input      [7:0]    io_write_payload,
  output              io_read_valid,
  input               io_read_ready,
  output     [7:0]    io_read_payload,
  output              io_uart_txd,
  input               io_uart_rxd,
  output              io_readError,
  input               io_writeBreak,
  output              io_readBreak,
  input               CLK_50,
  input               _zz_1
);
  wire                _zz_2;
  wire                tx_io_write_ready;
  wire                tx_io_txd;
  wire                rx_io_read_valid;
  wire       [7:0]    rx_io_read_payload;
  wire                rx_io_rts;
  wire                rx_io_error;
  wire                rx_io_break;
  reg        [19:0]   clockDivider_counter;
  wire                clockDivider_tick;
  reg                 io_write_thrown_valid;
  wire                io_write_thrown_ready;
  wire       [7:0]    io_write_thrown_payload;
  `ifndef SYNTHESIS
  reg [23:0] io_config_frame_stop_string;
  reg [31:0] io_config_frame_parity_string;
  `endif


  UartCtrlTx tx (
    .io_configFrame_dataLength    (io_config_frame_dataLength[2:0]  ), //i
    .io_configFrame_stop          (io_config_frame_stop             ), //i
    .io_configFrame_parity        (io_config_frame_parity[1:0]      ), //i
    .io_samplingTick              (clockDivider_tick                ), //i
    .io_write_valid               (io_write_thrown_valid            ), //i
    .io_write_ready               (tx_io_write_ready                ), //o
    .io_write_payload             (io_write_thrown_payload[7:0]     ), //i
    .io_cts                       (_zz_2                            ), //i
    .io_txd                       (tx_io_txd                        ), //o
    .io_break                     (io_writeBreak                    ), //i
    .CLK_50                       (CLK_50                           ), //i
    ._zz_2                        (_zz_1                            )  //i
  );
  UartCtrlRx rx (
    .io_configFrame_dataLength    (io_config_frame_dataLength[2:0]  ), //i
    .io_configFrame_stop          (io_config_frame_stop             ), //i
    .io_configFrame_parity        (io_config_frame_parity[1:0]      ), //i
    .io_samplingTick              (clockDivider_tick                ), //i
    .io_read_valid                (rx_io_read_valid                 ), //o
    .io_read_ready                (io_read_ready                    ), //i
    .io_read_payload              (rx_io_read_payload[7:0]          ), //o
    .io_rxd                       (io_uart_rxd                      ), //i
    .io_rts                       (rx_io_rts                        ), //o
    .io_error                     (rx_io_error                      ), //o
    .io_break                     (rx_io_break                      ), //o
    .CLK_50                       (CLK_50                           ), //i
    ._zz_2                        (_zz_1                            )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_config_frame_stop)
      `UartStopType_defaultEncoding_ONE : io_config_frame_stop_string = "ONE";
      `UartStopType_defaultEncoding_TWO : io_config_frame_stop_string = "TWO";
      default : io_config_frame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_config_frame_parity)
      `UartParityType_defaultEncoding_NONE : io_config_frame_parity_string = "NONE";
      `UartParityType_defaultEncoding_EVEN : io_config_frame_parity_string = "EVEN";
      `UartParityType_defaultEncoding_ODD : io_config_frame_parity_string = "ODD ";
      default : io_config_frame_parity_string = "????";
    endcase
  end
  `endif

  assign clockDivider_tick = (clockDivider_counter == 20'h0);
  always @ (*) begin
    io_write_thrown_valid = io_write_valid;
    if(rx_io_break)begin
      io_write_thrown_valid = 1'b0;
    end
  end

  always @ (*) begin
    io_write_ready = io_write_thrown_ready;
    if(rx_io_break)begin
      io_write_ready = 1'b1;
    end
  end

  assign io_write_thrown_payload = io_write_payload;
  assign io_write_thrown_ready = tx_io_write_ready;
  assign io_read_valid = rx_io_read_valid;
  assign io_read_payload = rx_io_read_payload;
  assign io_uart_txd = tx_io_txd;
  assign io_readError = rx_io_error;
  assign _zz_2 = 1'b0;
  assign io_readBreak = rx_io_break;
  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      clockDivider_counter <= 20'h0;
    end else begin
      clockDivider_counter <= (clockDivider_counter - 20'h00001);
      if(clockDivider_tick)begin
        clockDivider_counter <= io_config_clockDivider;
      end
    end
  end


endmodule

//UartCtrlRx replaced by UartCtrlRx

//UartCtrlTx replaced by UartCtrlTx

module Debounce (
  input      [102:0]  key_down,
  output              keyStatus_0_valid,
  output              keyStatus_0_payload,
  output              keyStatus_1_valid,
  output              keyStatus_1_payload,
  output              keyStatus_2_valid,
  output              keyStatus_2_payload,
  output              keyStatus_3_valid,
  output              keyStatus_3_payload,
  output              keyStatus_4_valid,
  output              keyStatus_4_payload,
  output              keyStatus_5_valid,
  output              keyStatus_5_payload,
  output              keyStatus_6_valid,
  output              keyStatus_6_payload,
  output              keyStatus_7_valid,
  output              keyStatus_7_payload,
  output              keyStatus_8_valid,
  output              keyStatus_8_payload,
  output              keyStatus_9_valid,
  output              keyStatus_9_payload,
  output              keyStatus_10_valid,
  output              keyStatus_10_payload,
  output              keyStatus_11_valid,
  output              keyStatus_11_payload,
  output              keyStatus_12_valid,
  output              keyStatus_12_payload,
  output              keyStatus_13_valid,
  output              keyStatus_13_payload,
  output              keyStatus_14_valid,
  output              keyStatus_14_payload,
  output              keyStatus_15_valid,
  output              keyStatus_15_payload,
  output              keyStatus_16_valid,
  output              keyStatus_16_payload,
  output              keyStatus_17_valid,
  output              keyStatus_17_payload,
  output              keyStatus_18_valid,
  output              keyStatus_18_payload,
  output              keyStatus_19_valid,
  output              keyStatus_19_payload,
  output              keyStatus_20_valid,
  output              keyStatus_20_payload,
  output              keyStatus_21_valid,
  output              keyStatus_21_payload,
  output              keyStatus_22_valid,
  output              keyStatus_22_payload,
  output              keyStatus_23_valid,
  output              keyStatus_23_payload,
  output              keyStatus_24_valid,
  output              keyStatus_24_payload,
  output              keyStatus_25_valid,
  output              keyStatus_25_payload,
  output              keyStatus_26_valid,
  output              keyStatus_26_payload,
  output              keyStatus_27_valid,
  output              keyStatus_27_payload,
  output              keyStatus_28_valid,
  output              keyStatus_28_payload,
  output              keyStatus_29_valid,
  output              keyStatus_29_payload,
  output              keyStatus_30_valid,
  output              keyStatus_30_payload,
  output              keyStatus_31_valid,
  output              keyStatus_31_payload,
  output              keyStatus_32_valid,
  output              keyStatus_32_payload,
  output              keyStatus_33_valid,
  output              keyStatus_33_payload,
  output              keyStatus_34_valid,
  output              keyStatus_34_payload,
  output              keyStatus_35_valid,
  output              keyStatus_35_payload,
  output              keyStatus_36_valid,
  output              keyStatus_36_payload,
  output              keyStatus_37_valid,
  output              keyStatus_37_payload,
  output              keyStatus_38_valid,
  output              keyStatus_38_payload,
  output              keyStatus_39_valid,
  output              keyStatus_39_payload,
  output              keyStatus_40_valid,
  output              keyStatus_40_payload,
  output              keyStatus_41_valid,
  output              keyStatus_41_payload,
  output              keyStatus_42_valid,
  output              keyStatus_42_payload,
  output              keyStatus_43_valid,
  output              keyStatus_43_payload,
  output              keyStatus_44_valid,
  output              keyStatus_44_payload,
  output              keyStatus_45_valid,
  output              keyStatus_45_payload,
  output              keyStatus_46_valid,
  output              keyStatus_46_payload,
  output              keyStatus_47_valid,
  output              keyStatus_47_payload,
  output              keyStatus_48_valid,
  output              keyStatus_48_payload,
  output              keyStatus_49_valid,
  output              keyStatus_49_payload,
  output              keyStatus_50_valid,
  output              keyStatus_50_payload,
  output              keyStatus_51_valid,
  output              keyStatus_51_payload,
  output              keyStatus_52_valid,
  output              keyStatus_52_payload,
  output              keyStatus_53_valid,
  output              keyStatus_53_payload,
  output              keyStatus_54_valid,
  output              keyStatus_54_payload,
  output              keyStatus_55_valid,
  output              keyStatus_55_payload,
  output              keyStatus_56_valid,
  output              keyStatus_56_payload,
  output              keyStatus_57_valid,
  output              keyStatus_57_payload,
  output              keyStatus_58_valid,
  output              keyStatus_58_payload,
  output              keyStatus_59_valid,
  output              keyStatus_59_payload,
  output              keyStatus_60_valid,
  output              keyStatus_60_payload,
  output              keyStatus_61_valid,
  output              keyStatus_61_payload,
  output              keyStatus_62_valid,
  output              keyStatus_62_payload,
  output              keyStatus_63_valid,
  output              keyStatus_63_payload,
  output              keyStatus_64_valid,
  output              keyStatus_64_payload,
  output              keyStatus_65_valid,
  output              keyStatus_65_payload,
  output              keyStatus_66_valid,
  output              keyStatus_66_payload,
  output              keyStatus_67_valid,
  output              keyStatus_67_payload,
  output              keyStatus_68_valid,
  output              keyStatus_68_payload,
  output              keyStatus_69_valid,
  output              keyStatus_69_payload,
  output              keyStatus_70_valid,
  output              keyStatus_70_payload,
  output              keyStatus_71_valid,
  output              keyStatus_71_payload,
  output              keyStatus_72_valid,
  output              keyStatus_72_payload,
  output              keyStatus_73_valid,
  output              keyStatus_73_payload,
  output              keyStatus_74_valid,
  output              keyStatus_74_payload,
  output              keyStatus_75_valid,
  output              keyStatus_75_payload,
  output              keyStatus_76_valid,
  output              keyStatus_76_payload,
  output              keyStatus_77_valid,
  output              keyStatus_77_payload,
  output              keyStatus_78_valid,
  output              keyStatus_78_payload,
  output              keyStatus_79_valid,
  output              keyStatus_79_payload,
  output              keyStatus_80_valid,
  output              keyStatus_80_payload,
  output              keyStatus_81_valid,
  output              keyStatus_81_payload,
  output              keyStatus_82_valid,
  output              keyStatus_82_payload,
  output              keyStatus_83_valid,
  output              keyStatus_83_payload,
  output              keyStatus_84_valid,
  output              keyStatus_84_payload,
  output              keyStatus_85_valid,
  output              keyStatus_85_payload,
  output              keyStatus_86_valid,
  output              keyStatus_86_payload,
  output              keyStatus_87_valid,
  output              keyStatus_87_payload,
  output              keyStatus_88_valid,
  output              keyStatus_88_payload,
  output              keyStatus_89_valid,
  output              keyStatus_89_payload,
  output              keyStatus_90_valid,
  output              keyStatus_90_payload,
  output              keyStatus_91_valid,
  output              keyStatus_91_payload,
  output              keyStatus_92_valid,
  output              keyStatus_92_payload,
  output              keyStatus_93_valid,
  output              keyStatus_93_payload,
  output              keyStatus_94_valid,
  output              keyStatus_94_payload,
  output              keyStatus_95_valid,
  output              keyStatus_95_payload,
  output              keyStatus_96_valid,
  output              keyStatus_96_payload,
  output              keyStatus_97_valid,
  output              keyStatus_97_payload,
  output              keyStatus_98_valid,
  output              keyStatus_98_payload,
  output              keyStatus_99_valid,
  output              keyStatus_99_payload,
  output              keyStatus_100_valid,
  output              keyStatus_100_payload,
  output              keyStatus_101_valid,
  output              keyStatus_101_payload,
  output              keyStatus_102_valid,
  output              keyStatus_102_payload,
  input               CLK_50,
  input               _zz_3
);
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                singleKey_103_filtered_valid;
  wire                singleKey_103_filtered_payload;
  wire                singleKey_104_filtered_valid;
  wire                singleKey_104_filtered_payload;
  wire                singleKey_105_filtered_valid;
  wire                singleKey_105_filtered_payload;
  wire                singleKey_106_filtered_valid;
  wire                singleKey_106_filtered_payload;
  wire                singleKey_107_filtered_valid;
  wire                singleKey_107_filtered_payload;
  wire                singleKey_108_filtered_valid;
  wire                singleKey_108_filtered_payload;
  wire                singleKey_109_filtered_valid;
  wire                singleKey_109_filtered_payload;
  wire                singleKey_110_filtered_valid;
  wire                singleKey_110_filtered_payload;
  wire                singleKey_111_filtered_valid;
  wire                singleKey_111_filtered_payload;
  wire                singleKey_112_filtered_valid;
  wire                singleKey_112_filtered_payload;
  wire                singleKey_113_filtered_valid;
  wire                singleKey_113_filtered_payload;
  wire                singleKey_114_filtered_valid;
  wire                singleKey_114_filtered_payload;
  wire                singleKey_115_filtered_valid;
  wire                singleKey_115_filtered_payload;
  wire                singleKey_116_filtered_valid;
  wire                singleKey_116_filtered_payload;
  wire                singleKey_117_filtered_valid;
  wire                singleKey_117_filtered_payload;
  wire                singleKey_118_filtered_valid;
  wire                singleKey_118_filtered_payload;
  wire                singleKey_119_filtered_valid;
  wire                singleKey_119_filtered_payload;
  wire                singleKey_120_filtered_valid;
  wire                singleKey_120_filtered_payload;
  wire                singleKey_121_filtered_valid;
  wire                singleKey_121_filtered_payload;
  wire                singleKey_122_filtered_valid;
  wire                singleKey_122_filtered_payload;
  wire                singleKey_123_filtered_valid;
  wire                singleKey_123_filtered_payload;
  wire                singleKey_124_filtered_valid;
  wire                singleKey_124_filtered_payload;
  wire                singleKey_125_filtered_valid;
  wire                singleKey_125_filtered_payload;
  wire                singleKey_126_filtered_valid;
  wire                singleKey_126_filtered_payload;
  wire                singleKey_127_filtered_valid;
  wire                singleKey_127_filtered_payload;
  wire                singleKey_128_filtered_valid;
  wire                singleKey_128_filtered_payload;
  wire                singleKey_129_filtered_valid;
  wire                singleKey_129_filtered_payload;
  wire                singleKey_130_filtered_valid;
  wire                singleKey_130_filtered_payload;
  wire                singleKey_131_filtered_valid;
  wire                singleKey_131_filtered_payload;
  wire                singleKey_132_filtered_valid;
  wire                singleKey_132_filtered_payload;
  wire                singleKey_133_filtered_valid;
  wire                singleKey_133_filtered_payload;
  wire                singleKey_134_filtered_valid;
  wire                singleKey_134_filtered_payload;
  wire                singleKey_135_filtered_valid;
  wire                singleKey_135_filtered_payload;
  wire                singleKey_136_filtered_valid;
  wire                singleKey_136_filtered_payload;
  wire                singleKey_137_filtered_valid;
  wire                singleKey_137_filtered_payload;
  wire                singleKey_138_filtered_valid;
  wire                singleKey_138_filtered_payload;
  wire                singleKey_139_filtered_valid;
  wire                singleKey_139_filtered_payload;
  wire                singleKey_140_filtered_valid;
  wire                singleKey_140_filtered_payload;
  wire                singleKey_141_filtered_valid;
  wire                singleKey_141_filtered_payload;
  wire                singleKey_142_filtered_valid;
  wire                singleKey_142_filtered_payload;
  wire                singleKey_143_filtered_valid;
  wire                singleKey_143_filtered_payload;
  wire                singleKey_144_filtered_valid;
  wire                singleKey_144_filtered_payload;
  wire                singleKey_145_filtered_valid;
  wire                singleKey_145_filtered_payload;
  wire                singleKey_146_filtered_valid;
  wire                singleKey_146_filtered_payload;
  wire                singleKey_147_filtered_valid;
  wire                singleKey_147_filtered_payload;
  wire                singleKey_148_filtered_valid;
  wire                singleKey_148_filtered_payload;
  wire                singleKey_149_filtered_valid;
  wire                singleKey_149_filtered_payload;
  wire                singleKey_150_filtered_valid;
  wire                singleKey_150_filtered_payload;
  wire                singleKey_151_filtered_valid;
  wire                singleKey_151_filtered_payload;
  wire                singleKey_152_filtered_valid;
  wire                singleKey_152_filtered_payload;
  wire                singleKey_153_filtered_valid;
  wire                singleKey_153_filtered_payload;
  wire                singleKey_154_filtered_valid;
  wire                singleKey_154_filtered_payload;
  wire                singleKey_155_filtered_valid;
  wire                singleKey_155_filtered_payload;
  wire                singleKey_156_filtered_valid;
  wire                singleKey_156_filtered_payload;
  wire                singleKey_157_filtered_valid;
  wire                singleKey_157_filtered_payload;
  wire                singleKey_158_filtered_valid;
  wire                singleKey_158_filtered_payload;
  wire                singleKey_159_filtered_valid;
  wire                singleKey_159_filtered_payload;
  wire                singleKey_160_filtered_valid;
  wire                singleKey_160_filtered_payload;
  wire                singleKey_161_filtered_valid;
  wire                singleKey_161_filtered_payload;
  wire                singleKey_162_filtered_valid;
  wire                singleKey_162_filtered_payload;
  wire                singleKey_163_filtered_valid;
  wire                singleKey_163_filtered_payload;
  wire                singleKey_164_filtered_valid;
  wire                singleKey_164_filtered_payload;
  wire                singleKey_165_filtered_valid;
  wire                singleKey_165_filtered_payload;
  wire                singleKey_166_filtered_valid;
  wire                singleKey_166_filtered_payload;
  wire                singleKey_167_filtered_valid;
  wire                singleKey_167_filtered_payload;
  wire                singleKey_168_filtered_valid;
  wire                singleKey_168_filtered_payload;
  wire                singleKey_169_filtered_valid;
  wire                singleKey_169_filtered_payload;
  wire                singleKey_170_filtered_valid;
  wire                singleKey_170_filtered_payload;
  wire                singleKey_171_filtered_valid;
  wire                singleKey_171_filtered_payload;
  wire                singleKey_172_filtered_valid;
  wire                singleKey_172_filtered_payload;
  wire                singleKey_173_filtered_valid;
  wire                singleKey_173_filtered_payload;
  wire                singleKey_174_filtered_valid;
  wire                singleKey_174_filtered_payload;
  wire                singleKey_175_filtered_valid;
  wire                singleKey_175_filtered_payload;
  wire                singleKey_176_filtered_valid;
  wire                singleKey_176_filtered_payload;
  wire                singleKey_177_filtered_valid;
  wire                singleKey_177_filtered_payload;
  wire                singleKey_178_filtered_valid;
  wire                singleKey_178_filtered_payload;
  wire                singleKey_179_filtered_valid;
  wire                singleKey_179_filtered_payload;
  wire                singleKey_180_filtered_valid;
  wire                singleKey_180_filtered_payload;
  wire                singleKey_181_filtered_valid;
  wire                singleKey_181_filtered_payload;
  wire                singleKey_182_filtered_valid;
  wire                singleKey_182_filtered_payload;
  wire                singleKey_183_filtered_valid;
  wire                singleKey_183_filtered_payload;
  wire                singleKey_184_filtered_valid;
  wire                singleKey_184_filtered_payload;
  wire                singleKey_185_filtered_valid;
  wire                singleKey_185_filtered_payload;
  wire                singleKey_186_filtered_valid;
  wire                singleKey_186_filtered_payload;
  wire                singleKey_187_filtered_valid;
  wire                singleKey_187_filtered_payload;
  wire                singleKey_188_filtered_valid;
  wire                singleKey_188_filtered_payload;
  wire                singleKey_189_filtered_valid;
  wire                singleKey_189_filtered_payload;
  wire                singleKey_190_filtered_valid;
  wire                singleKey_190_filtered_payload;
  wire                singleKey_191_filtered_valid;
  wire                singleKey_191_filtered_payload;
  wire                singleKey_192_filtered_valid;
  wire                singleKey_192_filtered_payload;
  wire                singleKey_193_filtered_valid;
  wire                singleKey_193_filtered_payload;
  wire                singleKey_194_filtered_valid;
  wire                singleKey_194_filtered_payload;
  wire                singleKey_195_filtered_valid;
  wire                singleKey_195_filtered_payload;
  wire                singleKey_196_filtered_valid;
  wire                singleKey_196_filtered_payload;
  wire                singleKey_197_filtered_valid;
  wire                singleKey_197_filtered_payload;
  wire                singleKey_198_filtered_valid;
  wire                singleKey_198_filtered_payload;
  wire                singleKey_199_filtered_valid;
  wire                singleKey_199_filtered_payload;
  wire                singleKey_200_filtered_valid;
  wire                singleKey_200_filtered_payload;
  wire                singleKey_201_filtered_valid;
  wire                singleKey_201_filtered_payload;
  wire                singleKey_202_filtered_valid;
  wire                singleKey_202_filtered_payload;
  wire                singleKey_203_filtered_valid;
  wire                singleKey_203_filtered_payload;
  wire                singleKey_204_filtered_valid;
  wire                singleKey_204_filtered_payload;
  wire                singleKey_205_filtered_valid;
  wire                singleKey_205_filtered_payload;
  reg        [14:0]   _zz_1;
  wire                _zz_2;
  reg                 _zz_2_regNext;

  SingleKey singleKey_103 (
    .raw                 (_zz_4                           ), //i
    .filtered_valid      (singleKey_103_filtered_valid    ), //o
    .filtered_payload    (singleKey_103_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_104 (
    .raw                 (_zz_5                           ), //i
    .filtered_valid      (singleKey_104_filtered_valid    ), //o
    .filtered_payload    (singleKey_104_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_105 (
    .raw                 (_zz_6                           ), //i
    .filtered_valid      (singleKey_105_filtered_valid    ), //o
    .filtered_payload    (singleKey_105_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_106 (
    .raw                 (_zz_7                           ), //i
    .filtered_valid      (singleKey_106_filtered_valid    ), //o
    .filtered_payload    (singleKey_106_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_107 (
    .raw                 (_zz_8                           ), //i
    .filtered_valid      (singleKey_107_filtered_valid    ), //o
    .filtered_payload    (singleKey_107_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_108 (
    .raw                 (_zz_9                           ), //i
    .filtered_valid      (singleKey_108_filtered_valid    ), //o
    .filtered_payload    (singleKey_108_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_109 (
    .raw                 (_zz_10                          ), //i
    .filtered_valid      (singleKey_109_filtered_valid    ), //o
    .filtered_payload    (singleKey_109_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_110 (
    .raw                 (_zz_11                          ), //i
    .filtered_valid      (singleKey_110_filtered_valid    ), //o
    .filtered_payload    (singleKey_110_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_111 (
    .raw                 (_zz_12                          ), //i
    .filtered_valid      (singleKey_111_filtered_valid    ), //o
    .filtered_payload    (singleKey_111_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_112 (
    .raw                 (_zz_13                          ), //i
    .filtered_valid      (singleKey_112_filtered_valid    ), //o
    .filtered_payload    (singleKey_112_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_113 (
    .raw                 (_zz_14                          ), //i
    .filtered_valid      (singleKey_113_filtered_valid    ), //o
    .filtered_payload    (singleKey_113_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_114 (
    .raw                 (_zz_15                          ), //i
    .filtered_valid      (singleKey_114_filtered_valid    ), //o
    .filtered_payload    (singleKey_114_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_115 (
    .raw                 (_zz_16                          ), //i
    .filtered_valid      (singleKey_115_filtered_valid    ), //o
    .filtered_payload    (singleKey_115_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_116 (
    .raw                 (_zz_17                          ), //i
    .filtered_valid      (singleKey_116_filtered_valid    ), //o
    .filtered_payload    (singleKey_116_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_117 (
    .raw                 (_zz_18                          ), //i
    .filtered_valid      (singleKey_117_filtered_valid    ), //o
    .filtered_payload    (singleKey_117_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_118 (
    .raw                 (_zz_19                          ), //i
    .filtered_valid      (singleKey_118_filtered_valid    ), //o
    .filtered_payload    (singleKey_118_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_119 (
    .raw                 (_zz_20                          ), //i
    .filtered_valid      (singleKey_119_filtered_valid    ), //o
    .filtered_payload    (singleKey_119_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_120 (
    .raw                 (_zz_21                          ), //i
    .filtered_valid      (singleKey_120_filtered_valid    ), //o
    .filtered_payload    (singleKey_120_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_121 (
    .raw                 (_zz_22                          ), //i
    .filtered_valid      (singleKey_121_filtered_valid    ), //o
    .filtered_payload    (singleKey_121_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_122 (
    .raw                 (_zz_23                          ), //i
    .filtered_valid      (singleKey_122_filtered_valid    ), //o
    .filtered_payload    (singleKey_122_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_123 (
    .raw                 (_zz_24                          ), //i
    .filtered_valid      (singleKey_123_filtered_valid    ), //o
    .filtered_payload    (singleKey_123_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_124 (
    .raw                 (_zz_25                          ), //i
    .filtered_valid      (singleKey_124_filtered_valid    ), //o
    .filtered_payload    (singleKey_124_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_125 (
    .raw                 (_zz_26                          ), //i
    .filtered_valid      (singleKey_125_filtered_valid    ), //o
    .filtered_payload    (singleKey_125_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_126 (
    .raw                 (_zz_27                          ), //i
    .filtered_valid      (singleKey_126_filtered_valid    ), //o
    .filtered_payload    (singleKey_126_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_127 (
    .raw                 (_zz_28                          ), //i
    .filtered_valid      (singleKey_127_filtered_valid    ), //o
    .filtered_payload    (singleKey_127_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_128 (
    .raw                 (_zz_29                          ), //i
    .filtered_valid      (singleKey_128_filtered_valid    ), //o
    .filtered_payload    (singleKey_128_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_129 (
    .raw                 (_zz_30                          ), //i
    .filtered_valid      (singleKey_129_filtered_valid    ), //o
    .filtered_payload    (singleKey_129_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_130 (
    .raw                 (_zz_31                          ), //i
    .filtered_valid      (singleKey_130_filtered_valid    ), //o
    .filtered_payload    (singleKey_130_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_131 (
    .raw                 (_zz_32                          ), //i
    .filtered_valid      (singleKey_131_filtered_valid    ), //o
    .filtered_payload    (singleKey_131_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_132 (
    .raw                 (_zz_33                          ), //i
    .filtered_valid      (singleKey_132_filtered_valid    ), //o
    .filtered_payload    (singleKey_132_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_133 (
    .raw                 (_zz_34                          ), //i
    .filtered_valid      (singleKey_133_filtered_valid    ), //o
    .filtered_payload    (singleKey_133_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_134 (
    .raw                 (_zz_35                          ), //i
    .filtered_valid      (singleKey_134_filtered_valid    ), //o
    .filtered_payload    (singleKey_134_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_135 (
    .raw                 (_zz_36                          ), //i
    .filtered_valid      (singleKey_135_filtered_valid    ), //o
    .filtered_payload    (singleKey_135_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_136 (
    .raw                 (_zz_37                          ), //i
    .filtered_valid      (singleKey_136_filtered_valid    ), //o
    .filtered_payload    (singleKey_136_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_137 (
    .raw                 (_zz_38                          ), //i
    .filtered_valid      (singleKey_137_filtered_valid    ), //o
    .filtered_payload    (singleKey_137_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_138 (
    .raw                 (_zz_39                          ), //i
    .filtered_valid      (singleKey_138_filtered_valid    ), //o
    .filtered_payload    (singleKey_138_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_139 (
    .raw                 (_zz_40                          ), //i
    .filtered_valid      (singleKey_139_filtered_valid    ), //o
    .filtered_payload    (singleKey_139_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_140 (
    .raw                 (_zz_41                          ), //i
    .filtered_valid      (singleKey_140_filtered_valid    ), //o
    .filtered_payload    (singleKey_140_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_141 (
    .raw                 (_zz_42                          ), //i
    .filtered_valid      (singleKey_141_filtered_valid    ), //o
    .filtered_payload    (singleKey_141_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_142 (
    .raw                 (_zz_43                          ), //i
    .filtered_valid      (singleKey_142_filtered_valid    ), //o
    .filtered_payload    (singleKey_142_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_143 (
    .raw                 (_zz_44                          ), //i
    .filtered_valid      (singleKey_143_filtered_valid    ), //o
    .filtered_payload    (singleKey_143_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_144 (
    .raw                 (_zz_45                          ), //i
    .filtered_valid      (singleKey_144_filtered_valid    ), //o
    .filtered_payload    (singleKey_144_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_145 (
    .raw                 (_zz_46                          ), //i
    .filtered_valid      (singleKey_145_filtered_valid    ), //o
    .filtered_payload    (singleKey_145_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_146 (
    .raw                 (_zz_47                          ), //i
    .filtered_valid      (singleKey_146_filtered_valid    ), //o
    .filtered_payload    (singleKey_146_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_147 (
    .raw                 (_zz_48                          ), //i
    .filtered_valid      (singleKey_147_filtered_valid    ), //o
    .filtered_payload    (singleKey_147_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_148 (
    .raw                 (_zz_49                          ), //i
    .filtered_valid      (singleKey_148_filtered_valid    ), //o
    .filtered_payload    (singleKey_148_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_149 (
    .raw                 (_zz_50                          ), //i
    .filtered_valid      (singleKey_149_filtered_valid    ), //o
    .filtered_payload    (singleKey_149_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_150 (
    .raw                 (_zz_51                          ), //i
    .filtered_valid      (singleKey_150_filtered_valid    ), //o
    .filtered_payload    (singleKey_150_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_151 (
    .raw                 (_zz_52                          ), //i
    .filtered_valid      (singleKey_151_filtered_valid    ), //o
    .filtered_payload    (singleKey_151_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_152 (
    .raw                 (_zz_53                          ), //i
    .filtered_valid      (singleKey_152_filtered_valid    ), //o
    .filtered_payload    (singleKey_152_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_153 (
    .raw                 (_zz_54                          ), //i
    .filtered_valid      (singleKey_153_filtered_valid    ), //o
    .filtered_payload    (singleKey_153_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_154 (
    .raw                 (_zz_55                          ), //i
    .filtered_valid      (singleKey_154_filtered_valid    ), //o
    .filtered_payload    (singleKey_154_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_155 (
    .raw                 (_zz_56                          ), //i
    .filtered_valid      (singleKey_155_filtered_valid    ), //o
    .filtered_payload    (singleKey_155_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_156 (
    .raw                 (_zz_57                          ), //i
    .filtered_valid      (singleKey_156_filtered_valid    ), //o
    .filtered_payload    (singleKey_156_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_157 (
    .raw                 (_zz_58                          ), //i
    .filtered_valid      (singleKey_157_filtered_valid    ), //o
    .filtered_payload    (singleKey_157_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_158 (
    .raw                 (_zz_59                          ), //i
    .filtered_valid      (singleKey_158_filtered_valid    ), //o
    .filtered_payload    (singleKey_158_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_159 (
    .raw                 (_zz_60                          ), //i
    .filtered_valid      (singleKey_159_filtered_valid    ), //o
    .filtered_payload    (singleKey_159_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_160 (
    .raw                 (_zz_61                          ), //i
    .filtered_valid      (singleKey_160_filtered_valid    ), //o
    .filtered_payload    (singleKey_160_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_161 (
    .raw                 (_zz_62                          ), //i
    .filtered_valid      (singleKey_161_filtered_valid    ), //o
    .filtered_payload    (singleKey_161_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_162 (
    .raw                 (_zz_63                          ), //i
    .filtered_valid      (singleKey_162_filtered_valid    ), //o
    .filtered_payload    (singleKey_162_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_163 (
    .raw                 (_zz_64                          ), //i
    .filtered_valid      (singleKey_163_filtered_valid    ), //o
    .filtered_payload    (singleKey_163_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_164 (
    .raw                 (_zz_65                          ), //i
    .filtered_valid      (singleKey_164_filtered_valid    ), //o
    .filtered_payload    (singleKey_164_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_165 (
    .raw                 (_zz_66                          ), //i
    .filtered_valid      (singleKey_165_filtered_valid    ), //o
    .filtered_payload    (singleKey_165_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_166 (
    .raw                 (_zz_67                          ), //i
    .filtered_valid      (singleKey_166_filtered_valid    ), //o
    .filtered_payload    (singleKey_166_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_167 (
    .raw                 (_zz_68                          ), //i
    .filtered_valid      (singleKey_167_filtered_valid    ), //o
    .filtered_payload    (singleKey_167_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_168 (
    .raw                 (_zz_69                          ), //i
    .filtered_valid      (singleKey_168_filtered_valid    ), //o
    .filtered_payload    (singleKey_168_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_169 (
    .raw                 (_zz_70                          ), //i
    .filtered_valid      (singleKey_169_filtered_valid    ), //o
    .filtered_payload    (singleKey_169_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_170 (
    .raw                 (_zz_71                          ), //i
    .filtered_valid      (singleKey_170_filtered_valid    ), //o
    .filtered_payload    (singleKey_170_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_171 (
    .raw                 (_zz_72                          ), //i
    .filtered_valid      (singleKey_171_filtered_valid    ), //o
    .filtered_payload    (singleKey_171_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_172 (
    .raw                 (_zz_73                          ), //i
    .filtered_valid      (singleKey_172_filtered_valid    ), //o
    .filtered_payload    (singleKey_172_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_173 (
    .raw                 (_zz_74                          ), //i
    .filtered_valid      (singleKey_173_filtered_valid    ), //o
    .filtered_payload    (singleKey_173_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_174 (
    .raw                 (_zz_75                          ), //i
    .filtered_valid      (singleKey_174_filtered_valid    ), //o
    .filtered_payload    (singleKey_174_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_175 (
    .raw                 (_zz_76                          ), //i
    .filtered_valid      (singleKey_175_filtered_valid    ), //o
    .filtered_payload    (singleKey_175_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_176 (
    .raw                 (_zz_77                          ), //i
    .filtered_valid      (singleKey_176_filtered_valid    ), //o
    .filtered_payload    (singleKey_176_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_177 (
    .raw                 (_zz_78                          ), //i
    .filtered_valid      (singleKey_177_filtered_valid    ), //o
    .filtered_payload    (singleKey_177_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_178 (
    .raw                 (_zz_79                          ), //i
    .filtered_valid      (singleKey_178_filtered_valid    ), //o
    .filtered_payload    (singleKey_178_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_179 (
    .raw                 (_zz_80                          ), //i
    .filtered_valid      (singleKey_179_filtered_valid    ), //o
    .filtered_payload    (singleKey_179_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_180 (
    .raw                 (_zz_81                          ), //i
    .filtered_valid      (singleKey_180_filtered_valid    ), //o
    .filtered_payload    (singleKey_180_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_181 (
    .raw                 (_zz_82                          ), //i
    .filtered_valid      (singleKey_181_filtered_valid    ), //o
    .filtered_payload    (singleKey_181_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_182 (
    .raw                 (_zz_83                          ), //i
    .filtered_valid      (singleKey_182_filtered_valid    ), //o
    .filtered_payload    (singleKey_182_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_183 (
    .raw                 (_zz_84                          ), //i
    .filtered_valid      (singleKey_183_filtered_valid    ), //o
    .filtered_payload    (singleKey_183_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_184 (
    .raw                 (_zz_85                          ), //i
    .filtered_valid      (singleKey_184_filtered_valid    ), //o
    .filtered_payload    (singleKey_184_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_185 (
    .raw                 (_zz_86                          ), //i
    .filtered_valid      (singleKey_185_filtered_valid    ), //o
    .filtered_payload    (singleKey_185_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_186 (
    .raw                 (_zz_87                          ), //i
    .filtered_valid      (singleKey_186_filtered_valid    ), //o
    .filtered_payload    (singleKey_186_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_187 (
    .raw                 (_zz_88                          ), //i
    .filtered_valid      (singleKey_187_filtered_valid    ), //o
    .filtered_payload    (singleKey_187_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_188 (
    .raw                 (_zz_89                          ), //i
    .filtered_valid      (singleKey_188_filtered_valid    ), //o
    .filtered_payload    (singleKey_188_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_189 (
    .raw                 (_zz_90                          ), //i
    .filtered_valid      (singleKey_189_filtered_valid    ), //o
    .filtered_payload    (singleKey_189_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_190 (
    .raw                 (_zz_91                          ), //i
    .filtered_valid      (singleKey_190_filtered_valid    ), //o
    .filtered_payload    (singleKey_190_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_191 (
    .raw                 (_zz_92                          ), //i
    .filtered_valid      (singleKey_191_filtered_valid    ), //o
    .filtered_payload    (singleKey_191_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_192 (
    .raw                 (_zz_93                          ), //i
    .filtered_valid      (singleKey_192_filtered_valid    ), //o
    .filtered_payload    (singleKey_192_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_193 (
    .raw                 (_zz_94                          ), //i
    .filtered_valid      (singleKey_193_filtered_valid    ), //o
    .filtered_payload    (singleKey_193_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_194 (
    .raw                 (_zz_95                          ), //i
    .filtered_valid      (singleKey_194_filtered_valid    ), //o
    .filtered_payload    (singleKey_194_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_195 (
    .raw                 (_zz_96                          ), //i
    .filtered_valid      (singleKey_195_filtered_valid    ), //o
    .filtered_payload    (singleKey_195_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_196 (
    .raw                 (_zz_97                          ), //i
    .filtered_valid      (singleKey_196_filtered_valid    ), //o
    .filtered_payload    (singleKey_196_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_197 (
    .raw                 (_zz_98                          ), //i
    .filtered_valid      (singleKey_197_filtered_valid    ), //o
    .filtered_payload    (singleKey_197_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_198 (
    .raw                 (_zz_99                          ), //i
    .filtered_valid      (singleKey_198_filtered_valid    ), //o
    .filtered_payload    (singleKey_198_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_199 (
    .raw                 (_zz_100                         ), //i
    .filtered_valid      (singleKey_199_filtered_valid    ), //o
    .filtered_payload    (singleKey_199_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_200 (
    .raw                 (_zz_101                         ), //i
    .filtered_valid      (singleKey_200_filtered_valid    ), //o
    .filtered_payload    (singleKey_200_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_201 (
    .raw                 (_zz_102                         ), //i
    .filtered_valid      (singleKey_201_filtered_valid    ), //o
    .filtered_payload    (singleKey_201_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_202 (
    .raw                 (_zz_103                         ), //i
    .filtered_valid      (singleKey_202_filtered_valid    ), //o
    .filtered_payload    (singleKey_202_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_203 (
    .raw                 (_zz_104                         ), //i
    .filtered_valid      (singleKey_203_filtered_valid    ), //o
    .filtered_payload    (singleKey_203_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_204 (
    .raw                 (_zz_105                         ), //i
    .filtered_valid      (singleKey_204_filtered_valid    ), //o
    .filtered_payload    (singleKey_204_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  SingleKey singleKey_205 (
    .raw                 (_zz_106                         ), //i
    .filtered_valid      (singleKey_205_filtered_valid    ), //o
    .filtered_payload    (singleKey_205_filtered_payload  ), //o
    .CLK_50              (CLK_50                          ), //i
    ._zz_3               (_zz_3                           ), //i
    ._zz_4               (_zz_2_regNext                   )  //i
  );
  assign _zz_2 = (_zz_1 == 15'h61a7);
  assign _zz_4 = key_down[0];
  assign keyStatus_0_valid = singleKey_103_filtered_valid;
  assign keyStatus_0_payload = singleKey_103_filtered_payload;
  assign _zz_5 = key_down[1];
  assign keyStatus_1_valid = singleKey_104_filtered_valid;
  assign keyStatus_1_payload = singleKey_104_filtered_payload;
  assign _zz_6 = key_down[2];
  assign keyStatus_2_valid = singleKey_105_filtered_valid;
  assign keyStatus_2_payload = singleKey_105_filtered_payload;
  assign _zz_7 = key_down[3];
  assign keyStatus_3_valid = singleKey_106_filtered_valid;
  assign keyStatus_3_payload = singleKey_106_filtered_payload;
  assign _zz_8 = key_down[4];
  assign keyStatus_4_valid = singleKey_107_filtered_valid;
  assign keyStatus_4_payload = singleKey_107_filtered_payload;
  assign _zz_9 = key_down[5];
  assign keyStatus_5_valid = singleKey_108_filtered_valid;
  assign keyStatus_5_payload = singleKey_108_filtered_payload;
  assign _zz_10 = key_down[6];
  assign keyStatus_6_valid = singleKey_109_filtered_valid;
  assign keyStatus_6_payload = singleKey_109_filtered_payload;
  assign _zz_11 = key_down[7];
  assign keyStatus_7_valid = singleKey_110_filtered_valid;
  assign keyStatus_7_payload = singleKey_110_filtered_payload;
  assign _zz_12 = key_down[8];
  assign keyStatus_8_valid = singleKey_111_filtered_valid;
  assign keyStatus_8_payload = singleKey_111_filtered_payload;
  assign _zz_13 = key_down[9];
  assign keyStatus_9_valid = singleKey_112_filtered_valid;
  assign keyStatus_9_payload = singleKey_112_filtered_payload;
  assign _zz_14 = key_down[10];
  assign keyStatus_10_valid = singleKey_113_filtered_valid;
  assign keyStatus_10_payload = singleKey_113_filtered_payload;
  assign _zz_15 = key_down[11];
  assign keyStatus_11_valid = singleKey_114_filtered_valid;
  assign keyStatus_11_payload = singleKey_114_filtered_payload;
  assign _zz_16 = key_down[12];
  assign keyStatus_12_valid = singleKey_115_filtered_valid;
  assign keyStatus_12_payload = singleKey_115_filtered_payload;
  assign _zz_17 = key_down[13];
  assign keyStatus_13_valid = singleKey_116_filtered_valid;
  assign keyStatus_13_payload = singleKey_116_filtered_payload;
  assign _zz_18 = key_down[14];
  assign keyStatus_14_valid = singleKey_117_filtered_valid;
  assign keyStatus_14_payload = singleKey_117_filtered_payload;
  assign _zz_19 = key_down[15];
  assign keyStatus_15_valid = singleKey_118_filtered_valid;
  assign keyStatus_15_payload = singleKey_118_filtered_payload;
  assign _zz_20 = key_down[16];
  assign keyStatus_16_valid = singleKey_119_filtered_valid;
  assign keyStatus_16_payload = singleKey_119_filtered_payload;
  assign _zz_21 = key_down[17];
  assign keyStatus_17_valid = singleKey_120_filtered_valid;
  assign keyStatus_17_payload = singleKey_120_filtered_payload;
  assign _zz_22 = key_down[18];
  assign keyStatus_18_valid = singleKey_121_filtered_valid;
  assign keyStatus_18_payload = singleKey_121_filtered_payload;
  assign _zz_23 = key_down[19];
  assign keyStatus_19_valid = singleKey_122_filtered_valid;
  assign keyStatus_19_payload = singleKey_122_filtered_payload;
  assign _zz_24 = key_down[20];
  assign keyStatus_20_valid = singleKey_123_filtered_valid;
  assign keyStatus_20_payload = singleKey_123_filtered_payload;
  assign _zz_25 = key_down[21];
  assign keyStatus_21_valid = singleKey_124_filtered_valid;
  assign keyStatus_21_payload = singleKey_124_filtered_payload;
  assign _zz_26 = key_down[22];
  assign keyStatus_22_valid = singleKey_125_filtered_valid;
  assign keyStatus_22_payload = singleKey_125_filtered_payload;
  assign _zz_27 = key_down[23];
  assign keyStatus_23_valid = singleKey_126_filtered_valid;
  assign keyStatus_23_payload = singleKey_126_filtered_payload;
  assign _zz_28 = key_down[24];
  assign keyStatus_24_valid = singleKey_127_filtered_valid;
  assign keyStatus_24_payload = singleKey_127_filtered_payload;
  assign _zz_29 = key_down[25];
  assign keyStatus_25_valid = singleKey_128_filtered_valid;
  assign keyStatus_25_payload = singleKey_128_filtered_payload;
  assign _zz_30 = key_down[26];
  assign keyStatus_26_valid = singleKey_129_filtered_valid;
  assign keyStatus_26_payload = singleKey_129_filtered_payload;
  assign _zz_31 = key_down[27];
  assign keyStatus_27_valid = singleKey_130_filtered_valid;
  assign keyStatus_27_payload = singleKey_130_filtered_payload;
  assign _zz_32 = key_down[28];
  assign keyStatus_28_valid = singleKey_131_filtered_valid;
  assign keyStatus_28_payload = singleKey_131_filtered_payload;
  assign _zz_33 = key_down[29];
  assign keyStatus_29_valid = singleKey_132_filtered_valid;
  assign keyStatus_29_payload = singleKey_132_filtered_payload;
  assign _zz_34 = key_down[30];
  assign keyStatus_30_valid = singleKey_133_filtered_valid;
  assign keyStatus_30_payload = singleKey_133_filtered_payload;
  assign _zz_35 = key_down[31];
  assign keyStatus_31_valid = singleKey_134_filtered_valid;
  assign keyStatus_31_payload = singleKey_134_filtered_payload;
  assign _zz_36 = key_down[32];
  assign keyStatus_32_valid = singleKey_135_filtered_valid;
  assign keyStatus_32_payload = singleKey_135_filtered_payload;
  assign _zz_37 = key_down[33];
  assign keyStatus_33_valid = singleKey_136_filtered_valid;
  assign keyStatus_33_payload = singleKey_136_filtered_payload;
  assign _zz_38 = key_down[34];
  assign keyStatus_34_valid = singleKey_137_filtered_valid;
  assign keyStatus_34_payload = singleKey_137_filtered_payload;
  assign _zz_39 = key_down[35];
  assign keyStatus_35_valid = singleKey_138_filtered_valid;
  assign keyStatus_35_payload = singleKey_138_filtered_payload;
  assign _zz_40 = key_down[36];
  assign keyStatus_36_valid = singleKey_139_filtered_valid;
  assign keyStatus_36_payload = singleKey_139_filtered_payload;
  assign _zz_41 = key_down[37];
  assign keyStatus_37_valid = singleKey_140_filtered_valid;
  assign keyStatus_37_payload = singleKey_140_filtered_payload;
  assign _zz_42 = key_down[38];
  assign keyStatus_38_valid = singleKey_141_filtered_valid;
  assign keyStatus_38_payload = singleKey_141_filtered_payload;
  assign _zz_43 = key_down[39];
  assign keyStatus_39_valid = singleKey_142_filtered_valid;
  assign keyStatus_39_payload = singleKey_142_filtered_payload;
  assign _zz_44 = key_down[40];
  assign keyStatus_40_valid = singleKey_143_filtered_valid;
  assign keyStatus_40_payload = singleKey_143_filtered_payload;
  assign _zz_45 = key_down[41];
  assign keyStatus_41_valid = singleKey_144_filtered_valid;
  assign keyStatus_41_payload = singleKey_144_filtered_payload;
  assign _zz_46 = key_down[42];
  assign keyStatus_42_valid = singleKey_145_filtered_valid;
  assign keyStatus_42_payload = singleKey_145_filtered_payload;
  assign _zz_47 = key_down[43];
  assign keyStatus_43_valid = singleKey_146_filtered_valid;
  assign keyStatus_43_payload = singleKey_146_filtered_payload;
  assign _zz_48 = key_down[44];
  assign keyStatus_44_valid = singleKey_147_filtered_valid;
  assign keyStatus_44_payload = singleKey_147_filtered_payload;
  assign _zz_49 = key_down[45];
  assign keyStatus_45_valid = singleKey_148_filtered_valid;
  assign keyStatus_45_payload = singleKey_148_filtered_payload;
  assign _zz_50 = key_down[46];
  assign keyStatus_46_valid = singleKey_149_filtered_valid;
  assign keyStatus_46_payload = singleKey_149_filtered_payload;
  assign _zz_51 = key_down[47];
  assign keyStatus_47_valid = singleKey_150_filtered_valid;
  assign keyStatus_47_payload = singleKey_150_filtered_payload;
  assign _zz_52 = key_down[48];
  assign keyStatus_48_valid = singleKey_151_filtered_valid;
  assign keyStatus_48_payload = singleKey_151_filtered_payload;
  assign _zz_53 = key_down[49];
  assign keyStatus_49_valid = singleKey_152_filtered_valid;
  assign keyStatus_49_payload = singleKey_152_filtered_payload;
  assign _zz_54 = key_down[50];
  assign keyStatus_50_valid = singleKey_153_filtered_valid;
  assign keyStatus_50_payload = singleKey_153_filtered_payload;
  assign _zz_55 = key_down[51];
  assign keyStatus_51_valid = singleKey_154_filtered_valid;
  assign keyStatus_51_payload = singleKey_154_filtered_payload;
  assign _zz_56 = key_down[52];
  assign keyStatus_52_valid = singleKey_155_filtered_valid;
  assign keyStatus_52_payload = singleKey_155_filtered_payload;
  assign _zz_57 = key_down[53];
  assign keyStatus_53_valid = singleKey_156_filtered_valid;
  assign keyStatus_53_payload = singleKey_156_filtered_payload;
  assign _zz_58 = key_down[54];
  assign keyStatus_54_valid = singleKey_157_filtered_valid;
  assign keyStatus_54_payload = singleKey_157_filtered_payload;
  assign _zz_59 = key_down[55];
  assign keyStatus_55_valid = singleKey_158_filtered_valid;
  assign keyStatus_55_payload = singleKey_158_filtered_payload;
  assign _zz_60 = key_down[56];
  assign keyStatus_56_valid = singleKey_159_filtered_valid;
  assign keyStatus_56_payload = singleKey_159_filtered_payload;
  assign _zz_61 = key_down[57];
  assign keyStatus_57_valid = singleKey_160_filtered_valid;
  assign keyStatus_57_payload = singleKey_160_filtered_payload;
  assign _zz_62 = key_down[58];
  assign keyStatus_58_valid = singleKey_161_filtered_valid;
  assign keyStatus_58_payload = singleKey_161_filtered_payload;
  assign _zz_63 = key_down[59];
  assign keyStatus_59_valid = singleKey_162_filtered_valid;
  assign keyStatus_59_payload = singleKey_162_filtered_payload;
  assign _zz_64 = key_down[60];
  assign keyStatus_60_valid = singleKey_163_filtered_valid;
  assign keyStatus_60_payload = singleKey_163_filtered_payload;
  assign _zz_65 = key_down[61];
  assign keyStatus_61_valid = singleKey_164_filtered_valid;
  assign keyStatus_61_payload = singleKey_164_filtered_payload;
  assign _zz_66 = key_down[62];
  assign keyStatus_62_valid = singleKey_165_filtered_valid;
  assign keyStatus_62_payload = singleKey_165_filtered_payload;
  assign _zz_67 = key_down[63];
  assign keyStatus_63_valid = singleKey_166_filtered_valid;
  assign keyStatus_63_payload = singleKey_166_filtered_payload;
  assign _zz_68 = key_down[64];
  assign keyStatus_64_valid = singleKey_167_filtered_valid;
  assign keyStatus_64_payload = singleKey_167_filtered_payload;
  assign _zz_69 = key_down[65];
  assign keyStatus_65_valid = singleKey_168_filtered_valid;
  assign keyStatus_65_payload = singleKey_168_filtered_payload;
  assign _zz_70 = key_down[66];
  assign keyStatus_66_valid = singleKey_169_filtered_valid;
  assign keyStatus_66_payload = singleKey_169_filtered_payload;
  assign _zz_71 = key_down[67];
  assign keyStatus_67_valid = singleKey_170_filtered_valid;
  assign keyStatus_67_payload = singleKey_170_filtered_payload;
  assign _zz_72 = key_down[68];
  assign keyStatus_68_valid = singleKey_171_filtered_valid;
  assign keyStatus_68_payload = singleKey_171_filtered_payload;
  assign _zz_73 = key_down[69];
  assign keyStatus_69_valid = singleKey_172_filtered_valid;
  assign keyStatus_69_payload = singleKey_172_filtered_payload;
  assign _zz_74 = key_down[70];
  assign keyStatus_70_valid = singleKey_173_filtered_valid;
  assign keyStatus_70_payload = singleKey_173_filtered_payload;
  assign _zz_75 = key_down[71];
  assign keyStatus_71_valid = singleKey_174_filtered_valid;
  assign keyStatus_71_payload = singleKey_174_filtered_payload;
  assign _zz_76 = key_down[72];
  assign keyStatus_72_valid = singleKey_175_filtered_valid;
  assign keyStatus_72_payload = singleKey_175_filtered_payload;
  assign _zz_77 = key_down[73];
  assign keyStatus_73_valid = singleKey_176_filtered_valid;
  assign keyStatus_73_payload = singleKey_176_filtered_payload;
  assign _zz_78 = key_down[74];
  assign keyStatus_74_valid = singleKey_177_filtered_valid;
  assign keyStatus_74_payload = singleKey_177_filtered_payload;
  assign _zz_79 = key_down[75];
  assign keyStatus_75_valid = singleKey_178_filtered_valid;
  assign keyStatus_75_payload = singleKey_178_filtered_payload;
  assign _zz_80 = key_down[76];
  assign keyStatus_76_valid = singleKey_179_filtered_valid;
  assign keyStatus_76_payload = singleKey_179_filtered_payload;
  assign _zz_81 = key_down[77];
  assign keyStatus_77_valid = singleKey_180_filtered_valid;
  assign keyStatus_77_payload = singleKey_180_filtered_payload;
  assign _zz_82 = key_down[78];
  assign keyStatus_78_valid = singleKey_181_filtered_valid;
  assign keyStatus_78_payload = singleKey_181_filtered_payload;
  assign _zz_83 = key_down[79];
  assign keyStatus_79_valid = singleKey_182_filtered_valid;
  assign keyStatus_79_payload = singleKey_182_filtered_payload;
  assign _zz_84 = key_down[80];
  assign keyStatus_80_valid = singleKey_183_filtered_valid;
  assign keyStatus_80_payload = singleKey_183_filtered_payload;
  assign _zz_85 = key_down[81];
  assign keyStatus_81_valid = singleKey_184_filtered_valid;
  assign keyStatus_81_payload = singleKey_184_filtered_payload;
  assign _zz_86 = key_down[82];
  assign keyStatus_82_valid = singleKey_185_filtered_valid;
  assign keyStatus_82_payload = singleKey_185_filtered_payload;
  assign _zz_87 = key_down[83];
  assign keyStatus_83_valid = singleKey_186_filtered_valid;
  assign keyStatus_83_payload = singleKey_186_filtered_payload;
  assign _zz_88 = key_down[84];
  assign keyStatus_84_valid = singleKey_187_filtered_valid;
  assign keyStatus_84_payload = singleKey_187_filtered_payload;
  assign _zz_89 = key_down[85];
  assign keyStatus_85_valid = singleKey_188_filtered_valid;
  assign keyStatus_85_payload = singleKey_188_filtered_payload;
  assign _zz_90 = key_down[86];
  assign keyStatus_86_valid = singleKey_189_filtered_valid;
  assign keyStatus_86_payload = singleKey_189_filtered_payload;
  assign _zz_91 = key_down[87];
  assign keyStatus_87_valid = singleKey_190_filtered_valid;
  assign keyStatus_87_payload = singleKey_190_filtered_payload;
  assign _zz_92 = key_down[88];
  assign keyStatus_88_valid = singleKey_191_filtered_valid;
  assign keyStatus_88_payload = singleKey_191_filtered_payload;
  assign _zz_93 = key_down[89];
  assign keyStatus_89_valid = singleKey_192_filtered_valid;
  assign keyStatus_89_payload = singleKey_192_filtered_payload;
  assign _zz_94 = key_down[90];
  assign keyStatus_90_valid = singleKey_193_filtered_valid;
  assign keyStatus_90_payload = singleKey_193_filtered_payload;
  assign _zz_95 = key_down[91];
  assign keyStatus_91_valid = singleKey_194_filtered_valid;
  assign keyStatus_91_payload = singleKey_194_filtered_payload;
  assign _zz_96 = key_down[92];
  assign keyStatus_92_valid = singleKey_195_filtered_valid;
  assign keyStatus_92_payload = singleKey_195_filtered_payload;
  assign _zz_97 = key_down[93];
  assign keyStatus_93_valid = singleKey_196_filtered_valid;
  assign keyStatus_93_payload = singleKey_196_filtered_payload;
  assign _zz_98 = key_down[94];
  assign keyStatus_94_valid = singleKey_197_filtered_valid;
  assign keyStatus_94_payload = singleKey_197_filtered_payload;
  assign _zz_99 = key_down[95];
  assign keyStatus_95_valid = singleKey_198_filtered_valid;
  assign keyStatus_95_payload = singleKey_198_filtered_payload;
  assign _zz_100 = key_down[96];
  assign keyStatus_96_valid = singleKey_199_filtered_valid;
  assign keyStatus_96_payload = singleKey_199_filtered_payload;
  assign _zz_101 = key_down[97];
  assign keyStatus_97_valid = singleKey_200_filtered_valid;
  assign keyStatus_97_payload = singleKey_200_filtered_payload;
  assign _zz_102 = key_down[98];
  assign keyStatus_98_valid = singleKey_201_filtered_valid;
  assign keyStatus_98_payload = singleKey_201_filtered_payload;
  assign _zz_103 = key_down[99];
  assign keyStatus_99_valid = singleKey_202_filtered_valid;
  assign keyStatus_99_payload = singleKey_202_filtered_payload;
  assign _zz_104 = key_down[100];
  assign keyStatus_100_valid = singleKey_203_filtered_valid;
  assign keyStatus_100_payload = singleKey_203_filtered_payload;
  assign _zz_105 = key_down[101];
  assign keyStatus_101_valid = singleKey_204_filtered_valid;
  assign keyStatus_101_payload = singleKey_204_filtered_payload;
  assign _zz_106 = key_down[102];
  assign keyStatus_102_valid = singleKey_205_filtered_valid;
  assign keyStatus_102_payload = singleKey_205_filtered_payload;
  always @ (posedge CLK_50 or posedge _zz_3) begin
    if (_zz_3) begin
      _zz_1 <= 15'h0;
      _zz_2_regNext <= 1'b0;
    end else begin
      _zz_1 <= (_zz_1 + 15'h0001);
      if(_zz_2)begin
        _zz_1 <= 15'h0;
      end
      _zz_2_regNext <= _zz_2;
    end
  end


endmodule

module UartCtrlRx (
  input      [2:0]    io_configFrame_dataLength,
  input      `UartStopType_defaultEncoding_type io_configFrame_stop,
  input      `UartParityType_defaultEncoding_type io_configFrame_parity,
  input               io_samplingTick,
  output              io_read_valid,
  input               io_read_ready,
  output     [7:0]    io_read_payload,
  input               io_rxd,
  output              io_rts,
  output reg          io_error,
  output              io_break,
  input               CLK_50,
  input               _zz_2
);
  wire                io_rxd_buffercc_io_dataOut;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire       [0:0]    _zz_7;
  wire       [2:0]    _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  reg                 _zz_1;
  wire                sampler_synchroniser;
  wire                sampler_samples_0;
  reg                 sampler_samples_1;
  reg                 sampler_samples_2;
  reg                 sampler_samples_3;
  reg                 sampler_samples_4;
  reg                 sampler_value;
  reg                 sampler_tick;
  reg        [2:0]    bitTimer_counter;
  reg                 bitTimer_tick;
  reg        [2:0]    bitCounter_value;
  reg        [6:0]    break_counter;
  wire                break_valid;
  reg        `UartCtrlRxState_defaultEncoding_type stateMachine_state;
  reg                 stateMachine_parity;
  reg        [7:0]    stateMachine_shifter;
  reg                 stateMachine_validReg;
  `ifndef SYNTHESIS
  reg [23:0] io_configFrame_stop_string;
  reg [31:0] io_configFrame_parity_string;
  reg [47:0] stateMachine_state_string;
  `endif


  assign _zz_3 = (stateMachine_parity == sampler_value);
  assign _zz_4 = (! sampler_value);
  assign _zz_5 = ((sampler_tick && (! sampler_value)) && (! break_valid));
  assign _zz_6 = (bitCounter_value == io_configFrame_dataLength);
  assign _zz_7 = ((io_configFrame_stop == `UartStopType_defaultEncoding_ONE) ? 1'b0 : 1'b1);
  assign _zz_8 = {2'd0, _zz_7};
  assign _zz_9 = ((((1'b0 || ((_zz_14 && sampler_samples_1) && sampler_samples_2)) || (((_zz_15 && sampler_samples_0) && sampler_samples_1) && sampler_samples_3)) || (((1'b1 && sampler_samples_0) && sampler_samples_2) && sampler_samples_3)) || (((1'b1 && sampler_samples_1) && sampler_samples_2) && sampler_samples_3));
  assign _zz_10 = (((1'b1 && sampler_samples_0) && sampler_samples_1) && sampler_samples_4);
  assign _zz_11 = ((1'b1 && sampler_samples_0) && sampler_samples_2);
  assign _zz_12 = (1'b1 && sampler_samples_1);
  assign _zz_13 = 1'b1;
  assign _zz_14 = (1'b1 && sampler_samples_0);
  assign _zz_15 = 1'b1;
  BufferCC io_rxd_buffercc (
    .io_dataIn     (io_rxd                      ), //i
    .io_dataOut    (io_rxd_buffercc_io_dataOut  ), //o
    .CLK_50        (CLK_50                      ), //i
    ._zz_1         (_zz_2                       )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_configFrame_stop)
      `UartStopType_defaultEncoding_ONE : io_configFrame_stop_string = "ONE";
      `UartStopType_defaultEncoding_TWO : io_configFrame_stop_string = "TWO";
      default : io_configFrame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_configFrame_parity)
      `UartParityType_defaultEncoding_NONE : io_configFrame_parity_string = "NONE";
      `UartParityType_defaultEncoding_EVEN : io_configFrame_parity_string = "EVEN";
      `UartParityType_defaultEncoding_ODD : io_configFrame_parity_string = "ODD ";
      default : io_configFrame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(stateMachine_state)
      `UartCtrlRxState_defaultEncoding_IDLE : stateMachine_state_string = "IDLE  ";
      `UartCtrlRxState_defaultEncoding_START : stateMachine_state_string = "START ";
      `UartCtrlRxState_defaultEncoding_DATA : stateMachine_state_string = "DATA  ";
      `UartCtrlRxState_defaultEncoding_PARITY : stateMachine_state_string = "PARITY";
      `UartCtrlRxState_defaultEncoding_STOP : stateMachine_state_string = "STOP  ";
      default : stateMachine_state_string = "??????";
    endcase
  end
  `endif

  always @ (*) begin
    io_error = 1'b0;
    case(stateMachine_state)
      `UartCtrlRxState_defaultEncoding_IDLE : begin
      end
      `UartCtrlRxState_defaultEncoding_START : begin
      end
      `UartCtrlRxState_defaultEncoding_DATA : begin
      end
      `UartCtrlRxState_defaultEncoding_PARITY : begin
        if(bitTimer_tick)begin
          if(! _zz_3) begin
            io_error = 1'b1;
          end
        end
      end
      default : begin
        if(bitTimer_tick)begin
          if(_zz_4)begin
            io_error = 1'b1;
          end
        end
      end
    endcase
  end

  assign io_rts = _zz_1;
  assign sampler_synchroniser = io_rxd_buffercc_io_dataOut;
  assign sampler_samples_0 = sampler_synchroniser;
  always @ (*) begin
    bitTimer_tick = 1'b0;
    if(sampler_tick)begin
      if((bitTimer_counter == 3'b000))begin
        bitTimer_tick = 1'b1;
      end
    end
  end

  assign break_valid = (break_counter == 7'h68);
  assign io_break = break_valid;
  assign io_read_valid = stateMachine_validReg;
  assign io_read_payload = stateMachine_shifter;
  always @ (posedge CLK_50 or posedge _zz_2) begin
    if (_zz_2) begin
      _zz_1 <= 1'b0;
      sampler_samples_1 <= 1'b1;
      sampler_samples_2 <= 1'b1;
      sampler_samples_3 <= 1'b1;
      sampler_samples_4 <= 1'b1;
      sampler_value <= 1'b1;
      sampler_tick <= 1'b0;
      break_counter <= 7'h0;
      stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
      stateMachine_validReg <= 1'b0;
    end else begin
      _zz_1 <= (! io_read_ready);
      if(io_samplingTick)begin
        sampler_samples_1 <= sampler_samples_0;
      end
      if(io_samplingTick)begin
        sampler_samples_2 <= sampler_samples_1;
      end
      if(io_samplingTick)begin
        sampler_samples_3 <= sampler_samples_2;
      end
      if(io_samplingTick)begin
        sampler_samples_4 <= sampler_samples_3;
      end
      sampler_value <= ((((((_zz_9 || _zz_10) || (_zz_11 && sampler_samples_4)) || ((_zz_12 && sampler_samples_2) && sampler_samples_4)) || (((_zz_13 && sampler_samples_0) && sampler_samples_3) && sampler_samples_4)) || (((1'b1 && sampler_samples_1) && sampler_samples_3) && sampler_samples_4)) || (((1'b1 && sampler_samples_2) && sampler_samples_3) && sampler_samples_4));
      sampler_tick <= io_samplingTick;
      if(sampler_value)begin
        break_counter <= 7'h0;
      end else begin
        if((io_samplingTick && (! break_valid)))begin
          break_counter <= (break_counter + 7'h01);
        end
      end
      stateMachine_validReg <= 1'b0;
      case(stateMachine_state)
        `UartCtrlRxState_defaultEncoding_IDLE : begin
          if(_zz_5)begin
            stateMachine_state <= `UartCtrlRxState_defaultEncoding_START;
          end
        end
        `UartCtrlRxState_defaultEncoding_START : begin
          if(bitTimer_tick)begin
            stateMachine_state <= `UartCtrlRxState_defaultEncoding_DATA;
            if((sampler_value == 1'b1))begin
              stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
            end
          end
        end
        `UartCtrlRxState_defaultEncoding_DATA : begin
          if(bitTimer_tick)begin
            if(_zz_6)begin
              if((io_configFrame_parity == `UartParityType_defaultEncoding_NONE))begin
                stateMachine_state <= `UartCtrlRxState_defaultEncoding_STOP;
                stateMachine_validReg <= 1'b1;
              end else begin
                stateMachine_state <= `UartCtrlRxState_defaultEncoding_PARITY;
              end
            end
          end
        end
        `UartCtrlRxState_defaultEncoding_PARITY : begin
          if(bitTimer_tick)begin
            if(_zz_3)begin
              stateMachine_state <= `UartCtrlRxState_defaultEncoding_STOP;
              stateMachine_validReg <= 1'b1;
            end else begin
              stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
            end
          end
        end
        default : begin
          if(bitTimer_tick)begin
            if(_zz_4)begin
              stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
            end else begin
              if((bitCounter_value == _zz_8))begin
                stateMachine_state <= `UartCtrlRxState_defaultEncoding_IDLE;
              end
            end
          end
        end
      endcase
    end
  end

  always @ (posedge CLK_50) begin
    if(sampler_tick)begin
      bitTimer_counter <= (bitTimer_counter - 3'b001);
    end
    if(bitTimer_tick)begin
      bitCounter_value <= (bitCounter_value + 3'b001);
    end
    if(bitTimer_tick)begin
      stateMachine_parity <= (stateMachine_parity ^ sampler_value);
    end
    case(stateMachine_state)
      `UartCtrlRxState_defaultEncoding_IDLE : begin
        if(_zz_5)begin
          bitTimer_counter <= 3'b010;
        end
      end
      `UartCtrlRxState_defaultEncoding_START : begin
        if(bitTimer_tick)begin
          bitCounter_value <= 3'b000;
          stateMachine_parity <= (io_configFrame_parity == `UartParityType_defaultEncoding_ODD);
        end
      end
      `UartCtrlRxState_defaultEncoding_DATA : begin
        if(bitTimer_tick)begin
          stateMachine_shifter[bitCounter_value] <= sampler_value;
          if(_zz_6)begin
            bitCounter_value <= 3'b000;
          end
        end
      end
      `UartCtrlRxState_defaultEncoding_PARITY : begin
        if(bitTimer_tick)begin
          bitCounter_value <= 3'b000;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module UartCtrlTx (
  input      [2:0]    io_configFrame_dataLength,
  input      `UartStopType_defaultEncoding_type io_configFrame_stop,
  input      `UartParityType_defaultEncoding_type io_configFrame_parity,
  input               io_samplingTick,
  input               io_write_valid,
  output reg          io_write_ready,
  input      [7:0]    io_write_payload,
  input               io_cts,
  output              io_txd,
  input               io_break,
  input               CLK_50,
  input               _zz_2
);
  wire                _zz_3;
  wire       [0:0]    _zz_4;
  wire       [2:0]    _zz_5;
  wire       [0:0]    _zz_6;
  wire       [2:0]    _zz_7;
  reg                 clockDivider_counter_willIncrement;
  wire                clockDivider_counter_willClear;
  reg        [2:0]    clockDivider_counter_valueNext;
  reg        [2:0]    clockDivider_counter_value;
  wire                clockDivider_counter_willOverflowIfInc;
  wire                clockDivider_counter_willOverflow;
  reg        [2:0]    tickCounter_value;
  reg        `UartCtrlTxState_defaultEncoding_type stateMachine_state;
  reg                 stateMachine_parity;
  reg                 stateMachine_txd;
  reg                 _zz_1;
  `ifndef SYNTHESIS
  reg [23:0] io_configFrame_stop_string;
  reg [31:0] io_configFrame_parity_string;
  reg [47:0] stateMachine_state_string;
  `endif


  assign _zz_3 = (tickCounter_value == io_configFrame_dataLength);
  assign _zz_4 = clockDivider_counter_willIncrement;
  assign _zz_5 = {2'd0, _zz_4};
  assign _zz_6 = ((io_configFrame_stop == `UartStopType_defaultEncoding_ONE) ? 1'b0 : 1'b1);
  assign _zz_7 = {2'd0, _zz_6};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_configFrame_stop)
      `UartStopType_defaultEncoding_ONE : io_configFrame_stop_string = "ONE";
      `UartStopType_defaultEncoding_TWO : io_configFrame_stop_string = "TWO";
      default : io_configFrame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_configFrame_parity)
      `UartParityType_defaultEncoding_NONE : io_configFrame_parity_string = "NONE";
      `UartParityType_defaultEncoding_EVEN : io_configFrame_parity_string = "EVEN";
      `UartParityType_defaultEncoding_ODD : io_configFrame_parity_string = "ODD ";
      default : io_configFrame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(stateMachine_state)
      `UartCtrlTxState_defaultEncoding_IDLE : stateMachine_state_string = "IDLE  ";
      `UartCtrlTxState_defaultEncoding_START : stateMachine_state_string = "START ";
      `UartCtrlTxState_defaultEncoding_DATA : stateMachine_state_string = "DATA  ";
      `UartCtrlTxState_defaultEncoding_PARITY : stateMachine_state_string = "PARITY";
      `UartCtrlTxState_defaultEncoding_STOP : stateMachine_state_string = "STOP  ";
      default : stateMachine_state_string = "??????";
    endcase
  end
  `endif

  always @ (*) begin
    clockDivider_counter_willIncrement = 1'b0;
    if(io_samplingTick)begin
      clockDivider_counter_willIncrement = 1'b1;
    end
  end

  assign clockDivider_counter_willClear = 1'b0;
  assign clockDivider_counter_willOverflowIfInc = (clockDivider_counter_value == 3'b111);
  assign clockDivider_counter_willOverflow = (clockDivider_counter_willOverflowIfInc && clockDivider_counter_willIncrement);
  always @ (*) begin
    clockDivider_counter_valueNext = (clockDivider_counter_value + _zz_5);
    if(clockDivider_counter_willClear)begin
      clockDivider_counter_valueNext = 3'b000;
    end
  end

  always @ (*) begin
    stateMachine_txd = 1'b1;
    case(stateMachine_state)
      `UartCtrlTxState_defaultEncoding_IDLE : begin
      end
      `UartCtrlTxState_defaultEncoding_START : begin
        stateMachine_txd = 1'b0;
      end
      `UartCtrlTxState_defaultEncoding_DATA : begin
        stateMachine_txd = io_write_payload[tickCounter_value];
      end
      `UartCtrlTxState_defaultEncoding_PARITY : begin
        stateMachine_txd = stateMachine_parity;
      end
      default : begin
      end
    endcase
  end

  always @ (*) begin
    io_write_ready = io_break;
    case(stateMachine_state)
      `UartCtrlTxState_defaultEncoding_IDLE : begin
      end
      `UartCtrlTxState_defaultEncoding_START : begin
      end
      `UartCtrlTxState_defaultEncoding_DATA : begin
        if(clockDivider_counter_willOverflow)begin
          if(_zz_3)begin
            io_write_ready = 1'b1;
          end
        end
      end
      `UartCtrlTxState_defaultEncoding_PARITY : begin
      end
      default : begin
      end
    endcase
  end

  assign io_txd = _zz_1;
  always @ (posedge CLK_50 or posedge _zz_2) begin
    if (_zz_2) begin
      clockDivider_counter_value <= 3'b000;
      stateMachine_state <= `UartCtrlTxState_defaultEncoding_IDLE;
      _zz_1 <= 1'b1;
    end else begin
      clockDivider_counter_value <= clockDivider_counter_valueNext;
      case(stateMachine_state)
        `UartCtrlTxState_defaultEncoding_IDLE : begin
          if(((io_write_valid && (! io_cts)) && clockDivider_counter_willOverflow))begin
            stateMachine_state <= `UartCtrlTxState_defaultEncoding_START;
          end
        end
        `UartCtrlTxState_defaultEncoding_START : begin
          if(clockDivider_counter_willOverflow)begin
            stateMachine_state <= `UartCtrlTxState_defaultEncoding_DATA;
          end
        end
        `UartCtrlTxState_defaultEncoding_DATA : begin
          if(clockDivider_counter_willOverflow)begin
            if(_zz_3)begin
              if((io_configFrame_parity == `UartParityType_defaultEncoding_NONE))begin
                stateMachine_state <= `UartCtrlTxState_defaultEncoding_STOP;
              end else begin
                stateMachine_state <= `UartCtrlTxState_defaultEncoding_PARITY;
              end
            end
          end
        end
        `UartCtrlTxState_defaultEncoding_PARITY : begin
          if(clockDivider_counter_willOverflow)begin
            stateMachine_state <= `UartCtrlTxState_defaultEncoding_STOP;
          end
        end
        default : begin
          if(clockDivider_counter_willOverflow)begin
            if((tickCounter_value == _zz_7))begin
              stateMachine_state <= (io_write_valid ? `UartCtrlTxState_defaultEncoding_START : `UartCtrlTxState_defaultEncoding_IDLE);
            end
          end
        end
      endcase
      _zz_1 <= (stateMachine_txd && (! io_break));
    end
  end

  always @ (posedge CLK_50) begin
    if(clockDivider_counter_willOverflow)begin
      tickCounter_value <= (tickCounter_value + 3'b001);
    end
    if(clockDivider_counter_willOverflow)begin
      stateMachine_parity <= (stateMachine_parity ^ stateMachine_txd);
    end
    case(stateMachine_state)
      `UartCtrlTxState_defaultEncoding_IDLE : begin
      end
      `UartCtrlTxState_defaultEncoding_START : begin
        if(clockDivider_counter_willOverflow)begin
          stateMachine_parity <= (io_configFrame_parity == `UartParityType_defaultEncoding_ODD);
          tickCounter_value <= 3'b000;
        end
      end
      `UartCtrlTxState_defaultEncoding_DATA : begin
        if(clockDivider_counter_willOverflow)begin
          if(_zz_3)begin
            tickCounter_value <= 3'b000;
          end
        end
      end
      `UartCtrlTxState_defaultEncoding_PARITY : begin
        if(clockDivider_counter_willOverflow)begin
          tickCounter_value <= 3'b000;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

//BufferCC replaced by BufferCC

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

//SingleKey replaced by SingleKey

module SingleKey (
  input               raw,
  output              filtered_valid,
  output              filtered_payload,
  input               CLK_50,
  input               _zz_3,
  input               _zz_4
);
  reg        [1:0]    cnt;
  reg                 raw_regNext;
  reg                 _zz_1;
  reg                 _zz_2;

  assign filtered_valid = _zz_1;
  assign filtered_payload = _zz_2;
  always @ (posedge CLK_50 or posedge _zz_3) begin
    if (_zz_3) begin
      cnt <= 2'b11;
    end else begin
      if(_zz_4) begin
        if((raw ^ raw_regNext))begin
          cnt <= 2'b11;
        end
        if((cnt != 2'b00))begin
          cnt <= (cnt - 2'b01);
        end
      end
    end
  end

  always @ (posedge CLK_50) begin
    if(_zz_4) begin
      raw_regNext <= raw;
      _zz_1 <= (cnt == 2'b01);
      if((cnt == 2'b01))begin
        _zz_2 <= (! raw);
      end
    end
  end


endmodule

module BufferCC (
  input               io_dataIn,
  output              io_dataOut,
  input               CLK_50,
  input               _zz_1
);
  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @ (posedge CLK_50 or posedge _zz_1) begin
    if (_zz_1) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule
